// ::BitSerialMatrixMultiplyTinyIO
module BitSerialMatrixMultiplyTinyIO(
	input clk,
	input wire  start,
	input wire [31:0] value,
	output /*mux_wire*/ logic  finish,
	output /*mux_wire*/ logic [31:0] result
);

/*state*/ logic [9:0][31:0] stored_values;
initial stored_values[0] = 'x;
initial stored_values[1] = 'x;
initial stored_values[2] = 'x;
initial stored_values[3] = 'x;
initial stored_values[4] = 'x;
initial stored_values[5] = 'x;
initial stored_values[6] = 'x;
initial stored_values[7] = 'x;
initial stored_values[8] = 'x;
initial stored_values[9] = 'x;
/*state*/ logic [31:0] last_value_use_as_addr;
initial last_value_use_as_addr = 'x;
/*latency*/ logic [31:0] _last_value_use_as_addr_D1; always_ff @(posedge clk) begin _last_value_use_as_addr_D1 <= last_value_use_as_addr; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D2; always_ff @(posedge clk) begin _last_value_use_as_addr_D2 <= _last_value_use_as_addr_D1; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D3; always_ff @(posedge clk) begin _last_value_use_as_addr_D3 <= _last_value_use_as_addr_D2; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D4; always_ff @(posedge clk) begin _last_value_use_as_addr_D4 <= _last_value_use_as_addr_D3; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D5; always_ff @(posedge clk) begin _last_value_use_as_addr_D5 <= _last_value_use_as_addr_D4; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D6; always_ff @(posedge clk) begin _last_value_use_as_addr_D6 <= _last_value_use_as_addr_D5; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D7; always_ff @(posedge clk) begin _last_value_use_as_addr_D7 <= _last_value_use_as_addr_D6; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D8; always_ff @(posedge clk) begin _last_value_use_as_addr_D8 <= _last_value_use_as_addr_D7; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D9; always_ff @(posedge clk) begin _last_value_use_as_addr_D9 <= _last_value_use_as_addr_D8; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D10; always_ff @(posedge clk) begin _last_value_use_as_addr_D10 <= _last_value_use_as_addr_D9; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D11; always_ff @(posedge clk) begin _last_value_use_as_addr_D11 <= _last_value_use_as_addr_D10; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D12; always_ff @(posedge clk) begin _last_value_use_as_addr_D12 <= _last_value_use_as_addr_D11; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D13; always_ff @(posedge clk) begin _last_value_use_as_addr_D13 <= _last_value_use_as_addr_D12; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D14; always_ff @(posedge clk) begin _last_value_use_as_addr_D14 <= _last_value_use_as_addr_D13; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D15; always_ff @(posedge clk) begin _last_value_use_as_addr_D15 <= _last_value_use_as_addr_D14; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D16; always_ff @(posedge clk) begin _last_value_use_as_addr_D16 <= _last_value_use_as_addr_D15; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D17; always_ff @(posedge clk) begin _last_value_use_as_addr_D17 <= _last_value_use_as_addr_D16; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D18; always_ff @(posedge clk) begin _last_value_use_as_addr_D18 <= _last_value_use_as_addr_D17; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D19; always_ff @(posedge clk) begin _last_value_use_as_addr_D19 <= _last_value_use_as_addr_D18; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D20; always_ff @(posedge clk) begin _last_value_use_as_addr_D20 <= _last_value_use_as_addr_D19; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D21; always_ff @(posedge clk) begin _last_value_use_as_addr_D21 <= _last_value_use_as_addr_D20; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D22; always_ff @(posedge clk) begin _last_value_use_as_addr_D22 <= _last_value_use_as_addr_D21; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D23; always_ff @(posedge clk) begin _last_value_use_as_addr_D23 <= _last_value_use_as_addr_D22; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D24; always_ff @(posedge clk) begin _last_value_use_as_addr_D24 <= _last_value_use_as_addr_D23; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D25; always_ff @(posedge clk) begin _last_value_use_as_addr_D25 <= _last_value_use_as_addr_D24; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D26; always_ff @(posedge clk) begin _last_value_use_as_addr_D26 <= _last_value_use_as_addr_D25; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D27; always_ff @(posedge clk) begin _last_value_use_as_addr_D27 <= _last_value_use_as_addr_D26; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D28; always_ff @(posedge clk) begin _last_value_use_as_addr_D28 <= _last_value_use_as_addr_D27; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D29; always_ff @(posedge clk) begin _last_value_use_as_addr_D29 <= _last_value_use_as_addr_D28; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D30; always_ff @(posedge clk) begin _last_value_use_as_addr_D30 <= _last_value_use_as_addr_D29; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D31; always_ff @(posedge clk) begin _last_value_use_as_addr_D31 <= _last_value_use_as_addr_D30; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D32; always_ff @(posedge clk) begin _last_value_use_as_addr_D32 <= _last_value_use_as_addr_D31; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D33; always_ff @(posedge clk) begin _last_value_use_as_addr_D33 <= _last_value_use_as_addr_D32; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D34; always_ff @(posedge clk) begin _last_value_use_as_addr_D34 <= _last_value_use_as_addr_D33; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D35; always_ff @(posedge clk) begin _last_value_use_as_addr_D35 <= _last_value_use_as_addr_D34; end
/*latency*/ logic [31:0] _last_value_use_as_addr_D36; always_ff @(posedge clk) begin _last_value_use_as_addr_D36 <= _last_value_use_as_addr_D35; end
/*mux_wire*/ logic [14:0][31:0] r;
/*mux_wire*/ logic  bsmm_start;
/*mux_wire*/ logic [9:0][31:0] bsmm_values;
wire  bsmm_finish;
wire [14:0][31:0] bsmm_result;
wire [31:0] _1 = r[_last_value_use_as_addr_D36];
BitSerialMatrixMultiplySpecific bsmm(
	.clk(clk),
	.start(bsmm_start),
	.values(bsmm_values),
	.finish(bsmm_finish),
	.result(bsmm_result)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	finish = 'x;
	finish = bsmm_finish;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	result = 'x;
	result = _1;
end
always_ff @(posedge clk) begin
	stored_values[last_value_use_as_addr] <= value;
end
always_ff @(posedge clk) begin
	last_value_use_as_addr <= value;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	r[0] = 'x;
	r[1] = 'x;
	r[2] = 'x;
	r[3] = 'x;
	r[4] = 'x;
	r[5] = 'x;
	r[6] = 'x;
	r[7] = 'x;
	r[8] = 'x;
	r[9] = 'x;
	r[10] = 'x;
	r[11] = 'x;
	r[12] = 'x;
	r[13] = 'x;
	r[14] = 'x;
	r = bsmm_result;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bsmm_start = 'x;
	bsmm_start = start;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bsmm_values[0] = 'x;
	bsmm_values[1] = 'x;
	bsmm_values[2] = 'x;
	bsmm_values[3] = 'x;
	bsmm_values[4] = 'x;
	bsmm_values[5] = 'x;
	bsmm_values[6] = 'x;
	bsmm_values[7] = 'x;
	bsmm_values[8] = 'x;
	bsmm_values[9] = 'x;
	bsmm_values = stored_values;
end
endmodule

// ::BitSerialMatrixMultiplySpecific
module BitSerialMatrixMultiplySpecific(
	input clk,
	input wire  start,
	input wire [9:0][31:0] values,
	output /*mux_wire*/ logic  finish,
	output /*mux_wire*/ logic [14:0][31:0] result
);

/*latency*/ logic  _start_D1; always_ff @(posedge clk) begin _start_D1 <= start; end
/*latency*/ logic  _start_D2; always_ff @(posedge clk) begin _start_D2 <= _start_D1; end
/*latency*/ logic  _start_D3; always_ff @(posedge clk) begin _start_D3 <= _start_D2; end
/*latency*/ logic  _start_D4; always_ff @(posedge clk) begin _start_D4 <= _start_D3; end
/*latency*/ logic  _start_D5; always_ff @(posedge clk) begin _start_D5 <= _start_D4; end
/*latency*/ logic  _start_D6; always_ff @(posedge clk) begin _start_D6 <= _start_D5; end
/*latency*/ logic  _start_D7; always_ff @(posedge clk) begin _start_D7 <= _start_D6; end
/*latency*/ logic  _start_D8; always_ff @(posedge clk) begin _start_D8 <= _start_D7; end
/*latency*/ logic  _start_D9; always_ff @(posedge clk) begin _start_D9 <= _start_D8; end
/*latency*/ logic  _start_D10; always_ff @(posedge clk) begin _start_D10 <= _start_D9; end
/*latency*/ logic  _start_D11; always_ff @(posedge clk) begin _start_D11 <= _start_D10; end
/*latency*/ logic  _start_D12; always_ff @(posedge clk) begin _start_D12 <= _start_D11; end
/*latency*/ logic  _start_D13; always_ff @(posedge clk) begin _start_D13 <= _start_D12; end
/*latency*/ logic  _start_D14; always_ff @(posedge clk) begin _start_D14 <= _start_D13; end
/*latency*/ logic  _start_D15; always_ff @(posedge clk) begin _start_D15 <= _start_D14; end
/*latency*/ logic  _start_D16; always_ff @(posedge clk) begin _start_D16 <= _start_D15; end
/*latency*/ logic  _start_D17; always_ff @(posedge clk) begin _start_D17 <= _start_D16; end
/*latency*/ logic  _start_D18; always_ff @(posedge clk) begin _start_D18 <= _start_D17; end
/*latency*/ logic  _start_D19; always_ff @(posedge clk) begin _start_D19 <= _start_D18; end
/*latency*/ logic  _start_D20; always_ff @(posedge clk) begin _start_D20 <= _start_D19; end
/*latency*/ logic  _start_D21; always_ff @(posedge clk) begin _start_D21 <= _start_D20; end
/*latency*/ logic  _start_D22; always_ff @(posedge clk) begin _start_D22 <= _start_D21; end
/*latency*/ logic  _start_D23; always_ff @(posedge clk) begin _start_D23 <= _start_D22; end
/*latency*/ logic  _start_D24; always_ff @(posedge clk) begin _start_D24 <= _start_D23; end
/*latency*/ logic  _start_D25; always_ff @(posedge clk) begin _start_D25 <= _start_D24; end
/*latency*/ logic  _start_D26; always_ff @(posedge clk) begin _start_D26 <= _start_D25; end
/*latency*/ logic  _start_D27; always_ff @(posedge clk) begin _start_D27 <= _start_D26; end
/*latency*/ logic  _start_D28; always_ff @(posedge clk) begin _start_D28 <= _start_D27; end
/*latency*/ logic  _start_D29; always_ff @(posedge clk) begin _start_D29 <= _start_D28; end
/*latency*/ logic  _start_D30; always_ff @(posedge clk) begin _start_D30 <= _start_D29; end
/*latency*/ logic  _start_D31; always_ff @(posedge clk) begin _start_D31 <= _start_D30; end
/*latency*/ logic  _start_D32; always_ff @(posedge clk) begin _start_D32 <= _start_D31; end
/*latency*/ logic  _start_D33; always_ff @(posedge clk) begin _start_D33 <= _start_D32; end
/*latency*/ logic  _start_D34; always_ff @(posedge clk) begin _start_D34 <= _start_D33; end
/*latency*/ logic  _start_D35; always_ff @(posedge clk) begin _start_D35 <= _start_D34; end
/*latency*/ logic  _start_D36; always_ff @(posedge clk) begin _start_D36 <= _start_D35; end
/*mux_wire*/ logic  bsmm_start;
/*mux_wire*/ logic [9:0][31:0] bsmm_values;
wire [14:0][31:0] bsmm_result;
BitSerialMatrixMultiply_WIDTH_10_HEIGHT_15_MATRIX___0_2_0_0_0_10_0_0_0_18___0_3_0_0_0_0_0_0_0_19___2_4_0_0_10_0_14_0_0_20___0_5_7_9_0_0_15_0_0_21___0_6_0_0_0_0_0_0_0_22___0_7_0_0_0_15_0_0_0_23___6_8_0_12_14_16_0_0_0_24___0_9_0_0_0_0_0_21_0_25___0_10_12_0_0_0_0_22_0_26___0_11_0_0_0_0_0_23_0_27___10_12_14_0_18_0_0_24_0_28___0_13_0_17_0_21_23_0_0_29___0_14_0_0_0_22_24_0_0_30___0_15_0_0_0_0_0_0_0_31___14_16_0_20_22_0_0_0_0_32___ bsmm(
	.clk(clk),
	.start(bsmm_start),
	.values(bsmm_values),
	.result(bsmm_result)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	finish = 'x;
	finish = _start_D36;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	result[0] = 'x;
	result[1] = 'x;
	result[2] = 'x;
	result[3] = 'x;
	result[4] = 'x;
	result[5] = 'x;
	result[6] = 'x;
	result[7] = 'x;
	result[8] = 'x;
	result[9] = 'x;
	result[10] = 'x;
	result[11] = 'x;
	result[12] = 'x;
	result[13] = 'x;
	result[14] = 'x;
	result = bsmm_result;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bsmm_start = 'x;
	bsmm_start = start;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bsmm_values[0] = 'x;
	bsmm_values[1] = 'x;
	bsmm_values[2] = 'x;
	bsmm_values[3] = 'x;
	bsmm_values[4] = 'x;
	bsmm_values[5] = 'x;
	bsmm_values[6] = 'x;
	bsmm_values[7] = 'x;
	bsmm_values[8] = 'x;
	bsmm_values[9] = 'x;
	bsmm_values = values;
end
endmodule

// ::BitSerialMatrixMultiply::<WIDTH = 10, HEIGHT = 15, MATRIX = [[0, 2, 0, 0, 0, 10, 0, 0, 0, 18], [0, 3, 0, 0, 0, 0, 0, 0, 0, 19], [2, 4, 0, 0, 10, 0, 14, 0, 0, 20], [0, 5, 7, 9, 0, 0, 15, 0, 0, 21], [0, 6, 0, 0, 0, 0, 0, 0, 0, 22], [0, 7, 0, 0, 0, 15, 0, 0, 0, 23], [6, 8, 0, 12, 14, 16, 0, 0, 0, 24], [0, 9, 0, 0, 0, 0, 0, 21, 0, 25], [0, 10, 12, 0, 0, 0, 0, 22, 0, 26], [0, 11, 0, 0, 0, 0, 0, 23, 0, 27], [10, 12, 14, 0, 18, 0, 0, 24, 0, 28], [0, 13, 0, 17, 0, 21, 23, 0, 0, 29], [0, 14, 0, 0, 0, 22, 24, 0, 0, 30], [0, 15, 0, 0, 0, 0, 0, 0, 0, 31], [14, 16, 0, 20, 22, 0, 0, 0, 0, 32]]>
module BitSerialMatrixMultiply_WIDTH_10_HEIGHT_15_MATRIX___0_2_0_0_0_10_0_0_0_18___0_3_0_0_0_0_0_0_0_19___2_4_0_0_10_0_14_0_0_20___0_5_7_9_0_0_15_0_0_21___0_6_0_0_0_0_0_0_0_22___0_7_0_0_0_15_0_0_0_23___6_8_0_12_14_16_0_0_0_24___0_9_0_0_0_0_0_21_0_25___0_10_12_0_0_0_0_22_0_26___0_11_0_0_0_0_0_23_0_27___10_12_14_0_18_0_0_24_0_28___0_13_0_17_0_21_23_0_0_29___0_14_0_0_0_22_24_0_0_30___0_15_0_0_0_0_0_0_0_31___14_16_0_20_22_0_0_0_0_32___(
	input clk,
	input wire  start,
	input wire [9:0][31:0] values,
	output /*mux_wire*/ logic [14:0][31:0] result
);

/*latency*/ logic  _start_D1; always_ff @(posedge clk) begin _start_D1 <= start; end
/*latency*/ logic  _start_D2; always_ff @(posedge clk) begin _start_D2 <= _start_D1; end
/*latency*/ logic  _start_D3; always_ff @(posedge clk) begin _start_D3 <= _start_D2; end
/*mux_wire*/ logic  shifter_start;
/*mux_wire*/ logic [9:0][31:0] shifter_values;
/*mux_wire*/ logic  bsm_state_start;
/*mux_wire*/ logic  iter_start;
/*mux_wire*/ logic [9:0] bits;
wire  iter_valid;
/*mux_wire*/ logic  shifter_shift;
wire [9:0] shifter_bits;
/*mux_wire*/ logic  bsm_state_feed;
/*mux_wire*/ logic [9:0] bsm_state_vector_bits;
wire [14:0][31:0] bsm_state_result_vector;
/*mux_wire*/ logic [14:0][31:0] _1_in;
wire [14:0][31:0] _1_out;
BitShifter_WIDTH_10_INT_BITWIDTH_32_ shifter(
	.clk(clk),
	.start(shifter_start),
	.values(shifter_values),
	.shift(shifter_shift),
	.bits(shifter_bits)
);
BitSerialMatrixMultiplyState_WIDTH_10_HEIGHT_15_MATRIX___0_2_0_0_0_10_0_0_0_18___0_3_0_0_0_0_0_0_0_19___2_4_0_0_10_0_14_0_0_20___0_5_7_9_0_0_15_0_0_21___0_6_0_0_0_0_0_0_0_22___0_7_0_0_0_15_0_0_0_23___6_8_0_12_14_16_0_0_0_24___0_9_0_0_0_0_0_21_0_25___0_10_12_0_0_0_0_22_0_26___0_11_0_0_0_0_0_23_0_27___10_12_14_0_18_0_0_24_0_28___0_13_0_17_0_21_23_0_0_29___0_14_0_0_0_22_24_0_0_30___0_15_0_0_0_0_0_0_0_31___14_16_0_20_22_0_0_0_0_32___ bsm_state(
	.clk(clk),
	.start(bsm_state_start),
	.feed(bsm_state_feed),
	.vector_bits(bsm_state_vector_bits),
	.result_vector(bsm_state_result_vector)
);
FixedSizeIterator_UP_TO_32_ iter(
	.clk(clk),
	.valid(iter_valid),
	.value(),
	.last(),
	.start(iter_start)
);
LatencyOffset_T_int_15__OFFSET_33_ _1(
	.clk(clk),
	.in(_1_in),
	.out(_1_out)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	result[0] = 'x;
	result[1] = 'x;
	result[2] = 'x;
	result[3] = 'x;
	result[4] = 'x;
	result[5] = 'x;
	result[6] = 'x;
	result[7] = 'x;
	result[8] = 'x;
	result[9] = 'x;
	result[10] = 'x;
	result[11] = 'x;
	result[12] = 'x;
	result[13] = 'x;
	result[14] = 'x;
	result = _1_out;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	shifter_start = 'x;
	shifter_start = start;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	shifter_values[0] = 'x;
	shifter_values[1] = 'x;
	shifter_values[2] = 'x;
	shifter_values[3] = 'x;
	shifter_values[4] = 'x;
	shifter_values[5] = 'x;
	shifter_values[6] = 'x;
	shifter_values[7] = 'x;
	shifter_values[8] = 'x;
	shifter_values[9] = 'x;
	shifter_values = values;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bsm_state_start = 'x;
	bsm_state_start = _start_D3;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	iter_start = 'x;
	iter_start = start;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bits[0] = 'x;
	bits[1] = 'x;
	bits[2] = 'x;
	bits[3] = 'x;
	bits[4] = 'x;
	bits[5] = 'x;
	bits[6] = 'x;
	bits[7] = 'x;
	bits[8] = 'x;
	bits[9] = 'x;
	bits = shifter_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	shifter_shift = 'x;
	shifter_shift = iter_valid;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bsm_state_feed = 'x;
	bsm_state_feed = iter_valid;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bsm_state_vector_bits[0] = 'x;
	bsm_state_vector_bits[1] = 'x;
	bsm_state_vector_bits[2] = 'x;
	bsm_state_vector_bits[3] = 'x;
	bsm_state_vector_bits[4] = 'x;
	bsm_state_vector_bits[5] = 'x;
	bsm_state_vector_bits[6] = 'x;
	bsm_state_vector_bits[7] = 'x;
	bsm_state_vector_bits[8] = 'x;
	bsm_state_vector_bits[9] = 'x;
	bsm_state_vector_bits = bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1_in[0] = 'x;
	_1_in[1] = 'x;
	_1_in[2] = 'x;
	_1_in[3] = 'x;
	_1_in[4] = 'x;
	_1_in[5] = 'x;
	_1_in[6] = 'x;
	_1_in[7] = 'x;
	_1_in[8] = 'x;
	_1_in[9] = 'x;
	_1_in[10] = 'x;
	_1_in[11] = 'x;
	_1_in[12] = 'x;
	_1_in[13] = 'x;
	_1_in[14] = 'x;
	_1_in = bsm_state_result_vector;
end
endmodule

// ::BitShifter::<WIDTH = 10, INT_BITWIDTH = 32>
module BitShifter_WIDTH_10_INT_BITWIDTH_32_(
	input clk,
	input wire  start,
	input wire [9:0][31:0] values,
	input wire  shift,
	output /*mux_wire*/ logic [9:0] bits
);

/*state*/ logic [31:0][9:0] split_into_bits;
initial split_into_bits[0][0] = 'x;
initial split_into_bits[0][1] = 'x;
initial split_into_bits[0][2] = 'x;
initial split_into_bits[0][3] = 'x;
initial split_into_bits[0][4] = 'x;
initial split_into_bits[0][5] = 'x;
initial split_into_bits[0][6] = 'x;
initial split_into_bits[0][7] = 'x;
initial split_into_bits[0][8] = 'x;
initial split_into_bits[0][9] = 'x;
initial split_into_bits[1][0] = 'x;
initial split_into_bits[1][1] = 'x;
initial split_into_bits[1][2] = 'x;
initial split_into_bits[1][3] = 'x;
initial split_into_bits[1][4] = 'x;
initial split_into_bits[1][5] = 'x;
initial split_into_bits[1][6] = 'x;
initial split_into_bits[1][7] = 'x;
initial split_into_bits[1][8] = 'x;
initial split_into_bits[1][9] = 'x;
initial split_into_bits[2][0] = 'x;
initial split_into_bits[2][1] = 'x;
initial split_into_bits[2][2] = 'x;
initial split_into_bits[2][3] = 'x;
initial split_into_bits[2][4] = 'x;
initial split_into_bits[2][5] = 'x;
initial split_into_bits[2][6] = 'x;
initial split_into_bits[2][7] = 'x;
initial split_into_bits[2][8] = 'x;
initial split_into_bits[2][9] = 'x;
initial split_into_bits[3][0] = 'x;
initial split_into_bits[3][1] = 'x;
initial split_into_bits[3][2] = 'x;
initial split_into_bits[3][3] = 'x;
initial split_into_bits[3][4] = 'x;
initial split_into_bits[3][5] = 'x;
initial split_into_bits[3][6] = 'x;
initial split_into_bits[3][7] = 'x;
initial split_into_bits[3][8] = 'x;
initial split_into_bits[3][9] = 'x;
initial split_into_bits[4][0] = 'x;
initial split_into_bits[4][1] = 'x;
initial split_into_bits[4][2] = 'x;
initial split_into_bits[4][3] = 'x;
initial split_into_bits[4][4] = 'x;
initial split_into_bits[4][5] = 'x;
initial split_into_bits[4][6] = 'x;
initial split_into_bits[4][7] = 'x;
initial split_into_bits[4][8] = 'x;
initial split_into_bits[4][9] = 'x;
initial split_into_bits[5][0] = 'x;
initial split_into_bits[5][1] = 'x;
initial split_into_bits[5][2] = 'x;
initial split_into_bits[5][3] = 'x;
initial split_into_bits[5][4] = 'x;
initial split_into_bits[5][5] = 'x;
initial split_into_bits[5][6] = 'x;
initial split_into_bits[5][7] = 'x;
initial split_into_bits[5][8] = 'x;
initial split_into_bits[5][9] = 'x;
initial split_into_bits[6][0] = 'x;
initial split_into_bits[6][1] = 'x;
initial split_into_bits[6][2] = 'x;
initial split_into_bits[6][3] = 'x;
initial split_into_bits[6][4] = 'x;
initial split_into_bits[6][5] = 'x;
initial split_into_bits[6][6] = 'x;
initial split_into_bits[6][7] = 'x;
initial split_into_bits[6][8] = 'x;
initial split_into_bits[6][9] = 'x;
initial split_into_bits[7][0] = 'x;
initial split_into_bits[7][1] = 'x;
initial split_into_bits[7][2] = 'x;
initial split_into_bits[7][3] = 'x;
initial split_into_bits[7][4] = 'x;
initial split_into_bits[7][5] = 'x;
initial split_into_bits[7][6] = 'x;
initial split_into_bits[7][7] = 'x;
initial split_into_bits[7][8] = 'x;
initial split_into_bits[7][9] = 'x;
initial split_into_bits[8][0] = 'x;
initial split_into_bits[8][1] = 'x;
initial split_into_bits[8][2] = 'x;
initial split_into_bits[8][3] = 'x;
initial split_into_bits[8][4] = 'x;
initial split_into_bits[8][5] = 'x;
initial split_into_bits[8][6] = 'x;
initial split_into_bits[8][7] = 'x;
initial split_into_bits[8][8] = 'x;
initial split_into_bits[8][9] = 'x;
initial split_into_bits[9][0] = 'x;
initial split_into_bits[9][1] = 'x;
initial split_into_bits[9][2] = 'x;
initial split_into_bits[9][3] = 'x;
initial split_into_bits[9][4] = 'x;
initial split_into_bits[9][5] = 'x;
initial split_into_bits[9][6] = 'x;
initial split_into_bits[9][7] = 'x;
initial split_into_bits[9][8] = 'x;
initial split_into_bits[9][9] = 'x;
initial split_into_bits[10][0] = 'x;
initial split_into_bits[10][1] = 'x;
initial split_into_bits[10][2] = 'x;
initial split_into_bits[10][3] = 'x;
initial split_into_bits[10][4] = 'x;
initial split_into_bits[10][5] = 'x;
initial split_into_bits[10][6] = 'x;
initial split_into_bits[10][7] = 'x;
initial split_into_bits[10][8] = 'x;
initial split_into_bits[10][9] = 'x;
initial split_into_bits[11][0] = 'x;
initial split_into_bits[11][1] = 'x;
initial split_into_bits[11][2] = 'x;
initial split_into_bits[11][3] = 'x;
initial split_into_bits[11][4] = 'x;
initial split_into_bits[11][5] = 'x;
initial split_into_bits[11][6] = 'x;
initial split_into_bits[11][7] = 'x;
initial split_into_bits[11][8] = 'x;
initial split_into_bits[11][9] = 'x;
initial split_into_bits[12][0] = 'x;
initial split_into_bits[12][1] = 'x;
initial split_into_bits[12][2] = 'x;
initial split_into_bits[12][3] = 'x;
initial split_into_bits[12][4] = 'x;
initial split_into_bits[12][5] = 'x;
initial split_into_bits[12][6] = 'x;
initial split_into_bits[12][7] = 'x;
initial split_into_bits[12][8] = 'x;
initial split_into_bits[12][9] = 'x;
initial split_into_bits[13][0] = 'x;
initial split_into_bits[13][1] = 'x;
initial split_into_bits[13][2] = 'x;
initial split_into_bits[13][3] = 'x;
initial split_into_bits[13][4] = 'x;
initial split_into_bits[13][5] = 'x;
initial split_into_bits[13][6] = 'x;
initial split_into_bits[13][7] = 'x;
initial split_into_bits[13][8] = 'x;
initial split_into_bits[13][9] = 'x;
initial split_into_bits[14][0] = 'x;
initial split_into_bits[14][1] = 'x;
initial split_into_bits[14][2] = 'x;
initial split_into_bits[14][3] = 'x;
initial split_into_bits[14][4] = 'x;
initial split_into_bits[14][5] = 'x;
initial split_into_bits[14][6] = 'x;
initial split_into_bits[14][7] = 'x;
initial split_into_bits[14][8] = 'x;
initial split_into_bits[14][9] = 'x;
initial split_into_bits[15][0] = 'x;
initial split_into_bits[15][1] = 'x;
initial split_into_bits[15][2] = 'x;
initial split_into_bits[15][3] = 'x;
initial split_into_bits[15][4] = 'x;
initial split_into_bits[15][5] = 'x;
initial split_into_bits[15][6] = 'x;
initial split_into_bits[15][7] = 'x;
initial split_into_bits[15][8] = 'x;
initial split_into_bits[15][9] = 'x;
initial split_into_bits[16][0] = 'x;
initial split_into_bits[16][1] = 'x;
initial split_into_bits[16][2] = 'x;
initial split_into_bits[16][3] = 'x;
initial split_into_bits[16][4] = 'x;
initial split_into_bits[16][5] = 'x;
initial split_into_bits[16][6] = 'x;
initial split_into_bits[16][7] = 'x;
initial split_into_bits[16][8] = 'x;
initial split_into_bits[16][9] = 'x;
initial split_into_bits[17][0] = 'x;
initial split_into_bits[17][1] = 'x;
initial split_into_bits[17][2] = 'x;
initial split_into_bits[17][3] = 'x;
initial split_into_bits[17][4] = 'x;
initial split_into_bits[17][5] = 'x;
initial split_into_bits[17][6] = 'x;
initial split_into_bits[17][7] = 'x;
initial split_into_bits[17][8] = 'x;
initial split_into_bits[17][9] = 'x;
initial split_into_bits[18][0] = 'x;
initial split_into_bits[18][1] = 'x;
initial split_into_bits[18][2] = 'x;
initial split_into_bits[18][3] = 'x;
initial split_into_bits[18][4] = 'x;
initial split_into_bits[18][5] = 'x;
initial split_into_bits[18][6] = 'x;
initial split_into_bits[18][7] = 'x;
initial split_into_bits[18][8] = 'x;
initial split_into_bits[18][9] = 'x;
initial split_into_bits[19][0] = 'x;
initial split_into_bits[19][1] = 'x;
initial split_into_bits[19][2] = 'x;
initial split_into_bits[19][3] = 'x;
initial split_into_bits[19][4] = 'x;
initial split_into_bits[19][5] = 'x;
initial split_into_bits[19][6] = 'x;
initial split_into_bits[19][7] = 'x;
initial split_into_bits[19][8] = 'x;
initial split_into_bits[19][9] = 'x;
initial split_into_bits[20][0] = 'x;
initial split_into_bits[20][1] = 'x;
initial split_into_bits[20][2] = 'x;
initial split_into_bits[20][3] = 'x;
initial split_into_bits[20][4] = 'x;
initial split_into_bits[20][5] = 'x;
initial split_into_bits[20][6] = 'x;
initial split_into_bits[20][7] = 'x;
initial split_into_bits[20][8] = 'x;
initial split_into_bits[20][9] = 'x;
initial split_into_bits[21][0] = 'x;
initial split_into_bits[21][1] = 'x;
initial split_into_bits[21][2] = 'x;
initial split_into_bits[21][3] = 'x;
initial split_into_bits[21][4] = 'x;
initial split_into_bits[21][5] = 'x;
initial split_into_bits[21][6] = 'x;
initial split_into_bits[21][7] = 'x;
initial split_into_bits[21][8] = 'x;
initial split_into_bits[21][9] = 'x;
initial split_into_bits[22][0] = 'x;
initial split_into_bits[22][1] = 'x;
initial split_into_bits[22][2] = 'x;
initial split_into_bits[22][3] = 'x;
initial split_into_bits[22][4] = 'x;
initial split_into_bits[22][5] = 'x;
initial split_into_bits[22][6] = 'x;
initial split_into_bits[22][7] = 'x;
initial split_into_bits[22][8] = 'x;
initial split_into_bits[22][9] = 'x;
initial split_into_bits[23][0] = 'x;
initial split_into_bits[23][1] = 'x;
initial split_into_bits[23][2] = 'x;
initial split_into_bits[23][3] = 'x;
initial split_into_bits[23][4] = 'x;
initial split_into_bits[23][5] = 'x;
initial split_into_bits[23][6] = 'x;
initial split_into_bits[23][7] = 'x;
initial split_into_bits[23][8] = 'x;
initial split_into_bits[23][9] = 'x;
initial split_into_bits[24][0] = 'x;
initial split_into_bits[24][1] = 'x;
initial split_into_bits[24][2] = 'x;
initial split_into_bits[24][3] = 'x;
initial split_into_bits[24][4] = 'x;
initial split_into_bits[24][5] = 'x;
initial split_into_bits[24][6] = 'x;
initial split_into_bits[24][7] = 'x;
initial split_into_bits[24][8] = 'x;
initial split_into_bits[24][9] = 'x;
initial split_into_bits[25][0] = 'x;
initial split_into_bits[25][1] = 'x;
initial split_into_bits[25][2] = 'x;
initial split_into_bits[25][3] = 'x;
initial split_into_bits[25][4] = 'x;
initial split_into_bits[25][5] = 'x;
initial split_into_bits[25][6] = 'x;
initial split_into_bits[25][7] = 'x;
initial split_into_bits[25][8] = 'x;
initial split_into_bits[25][9] = 'x;
initial split_into_bits[26][0] = 'x;
initial split_into_bits[26][1] = 'x;
initial split_into_bits[26][2] = 'x;
initial split_into_bits[26][3] = 'x;
initial split_into_bits[26][4] = 'x;
initial split_into_bits[26][5] = 'x;
initial split_into_bits[26][6] = 'x;
initial split_into_bits[26][7] = 'x;
initial split_into_bits[26][8] = 'x;
initial split_into_bits[26][9] = 'x;
initial split_into_bits[27][0] = 'x;
initial split_into_bits[27][1] = 'x;
initial split_into_bits[27][2] = 'x;
initial split_into_bits[27][3] = 'x;
initial split_into_bits[27][4] = 'x;
initial split_into_bits[27][5] = 'x;
initial split_into_bits[27][6] = 'x;
initial split_into_bits[27][7] = 'x;
initial split_into_bits[27][8] = 'x;
initial split_into_bits[27][9] = 'x;
initial split_into_bits[28][0] = 'x;
initial split_into_bits[28][1] = 'x;
initial split_into_bits[28][2] = 'x;
initial split_into_bits[28][3] = 'x;
initial split_into_bits[28][4] = 'x;
initial split_into_bits[28][5] = 'x;
initial split_into_bits[28][6] = 'x;
initial split_into_bits[28][7] = 'x;
initial split_into_bits[28][8] = 'x;
initial split_into_bits[28][9] = 'x;
initial split_into_bits[29][0] = 'x;
initial split_into_bits[29][1] = 'x;
initial split_into_bits[29][2] = 'x;
initial split_into_bits[29][3] = 'x;
initial split_into_bits[29][4] = 'x;
initial split_into_bits[29][5] = 'x;
initial split_into_bits[29][6] = 'x;
initial split_into_bits[29][7] = 'x;
initial split_into_bits[29][8] = 'x;
initial split_into_bits[29][9] = 'x;
initial split_into_bits[30][0] = 'x;
initial split_into_bits[30][1] = 'x;
initial split_into_bits[30][2] = 'x;
initial split_into_bits[30][3] = 'x;
initial split_into_bits[30][4] = 'x;
initial split_into_bits[30][5] = 'x;
initial split_into_bits[30][6] = 'x;
initial split_into_bits[30][7] = 'x;
initial split_into_bits[30][8] = 'x;
initial split_into_bits[30][9] = 'x;
initial split_into_bits[31][0] = 'x;
initial split_into_bits[31][1] = 'x;
initial split_into_bits[31][2] = 'x;
initial split_into_bits[31][3] = 'x;
initial split_into_bits[31][4] = 'x;
initial split_into_bits[31][5] = 'x;
initial split_into_bits[31][6] = 'x;
initial split_into_bits[31][7] = 'x;
initial split_into_bits[31][8] = 'x;
initial split_into_bits[31][9] = 'x;
/*mux_wire*/ logic [31:0] value_bits;
wire [31:0] _3 = values[0];
/*mux_wire*/ logic [31:0] _1_value;
wire [31:0] _1_bits;
wire  _5 = value_bits[0];
wire  _9 = value_bits[1];
wire  _13 = value_bits[2];
wire  _17 = value_bits[3];
wire  _21 = value_bits[4];
wire  _25 = value_bits[5];
wire  _29 = value_bits[6];
wire  _33 = value_bits[7];
wire  _37 = value_bits[8];
wire  _41 = value_bits[9];
wire  _45 = value_bits[10];
wire  _49 = value_bits[11];
wire  _53 = value_bits[12];
wire  _57 = value_bits[13];
wire  _61 = value_bits[14];
wire  _65 = value_bits[15];
wire  _69 = value_bits[16];
wire  _73 = value_bits[17];
wire  _77 = value_bits[18];
wire  _81 = value_bits[19];
wire  _85 = value_bits[20];
wire  _89 = value_bits[21];
wire  _93 = value_bits[22];
wire  _97 = value_bits[23];
wire  _101 = value_bits[24];
wire  _105 = value_bits[25];
wire  _109 = value_bits[26];
wire  _113 = value_bits[27];
wire  _117 = value_bits[28];
wire  _121 = value_bits[29];
wire  _125 = value_bits[30];
wire  _129 = value_bits[31];
/*mux_wire*/ logic [31:0] value_bits_2;
wire [31:0] _134 = values[1];
/*mux_wire*/ logic [31:0] _132_value;
wire [31:0] _132_bits;
wire  _136 = value_bits_2[0];
wire  _140 = value_bits_2[1];
wire  _144 = value_bits_2[2];
wire  _148 = value_bits_2[3];
wire  _152 = value_bits_2[4];
wire  _156 = value_bits_2[5];
wire  _160 = value_bits_2[6];
wire  _164 = value_bits_2[7];
wire  _168 = value_bits_2[8];
wire  _172 = value_bits_2[9];
wire  _176 = value_bits_2[10];
wire  _180 = value_bits_2[11];
wire  _184 = value_bits_2[12];
wire  _188 = value_bits_2[13];
wire  _192 = value_bits_2[14];
wire  _196 = value_bits_2[15];
wire  _200 = value_bits_2[16];
wire  _204 = value_bits_2[17];
wire  _208 = value_bits_2[18];
wire  _212 = value_bits_2[19];
wire  _216 = value_bits_2[20];
wire  _220 = value_bits_2[21];
wire  _224 = value_bits_2[22];
wire  _228 = value_bits_2[23];
wire  _232 = value_bits_2[24];
wire  _236 = value_bits_2[25];
wire  _240 = value_bits_2[26];
wire  _244 = value_bits_2[27];
wire  _248 = value_bits_2[28];
wire  _252 = value_bits_2[29];
wire  _256 = value_bits_2[30];
wire  _260 = value_bits_2[31];
/*mux_wire*/ logic [31:0] value_bits_3;
wire [31:0] _265 = values[2];
/*mux_wire*/ logic [31:0] _263_value;
wire [31:0] _263_bits;
wire  _267 = value_bits_3[0];
wire  _271 = value_bits_3[1];
wire  _275 = value_bits_3[2];
wire  _279 = value_bits_3[3];
wire  _283 = value_bits_3[4];
wire  _287 = value_bits_3[5];
wire  _291 = value_bits_3[6];
wire  _295 = value_bits_3[7];
wire  _299 = value_bits_3[8];
wire  _303 = value_bits_3[9];
wire  _307 = value_bits_3[10];
wire  _311 = value_bits_3[11];
wire  _315 = value_bits_3[12];
wire  _319 = value_bits_3[13];
wire  _323 = value_bits_3[14];
wire  _327 = value_bits_3[15];
wire  _331 = value_bits_3[16];
wire  _335 = value_bits_3[17];
wire  _339 = value_bits_3[18];
wire  _343 = value_bits_3[19];
wire  _347 = value_bits_3[20];
wire  _351 = value_bits_3[21];
wire  _355 = value_bits_3[22];
wire  _359 = value_bits_3[23];
wire  _363 = value_bits_3[24];
wire  _367 = value_bits_3[25];
wire  _371 = value_bits_3[26];
wire  _375 = value_bits_3[27];
wire  _379 = value_bits_3[28];
wire  _383 = value_bits_3[29];
wire  _387 = value_bits_3[30];
wire  _391 = value_bits_3[31];
/*mux_wire*/ logic [31:0] value_bits_4;
wire [31:0] _396 = values[3];
/*mux_wire*/ logic [31:0] _394_value;
wire [31:0] _394_bits;
wire  _398 = value_bits_4[0];
wire  _402 = value_bits_4[1];
wire  _406 = value_bits_4[2];
wire  _410 = value_bits_4[3];
wire  _414 = value_bits_4[4];
wire  _418 = value_bits_4[5];
wire  _422 = value_bits_4[6];
wire  _426 = value_bits_4[7];
wire  _430 = value_bits_4[8];
wire  _434 = value_bits_4[9];
wire  _438 = value_bits_4[10];
wire  _442 = value_bits_4[11];
wire  _446 = value_bits_4[12];
wire  _450 = value_bits_4[13];
wire  _454 = value_bits_4[14];
wire  _458 = value_bits_4[15];
wire  _462 = value_bits_4[16];
wire  _466 = value_bits_4[17];
wire  _470 = value_bits_4[18];
wire  _474 = value_bits_4[19];
wire  _478 = value_bits_4[20];
wire  _482 = value_bits_4[21];
wire  _486 = value_bits_4[22];
wire  _490 = value_bits_4[23];
wire  _494 = value_bits_4[24];
wire  _498 = value_bits_4[25];
wire  _502 = value_bits_4[26];
wire  _506 = value_bits_4[27];
wire  _510 = value_bits_4[28];
wire  _514 = value_bits_4[29];
wire  _518 = value_bits_4[30];
wire  _522 = value_bits_4[31];
/*mux_wire*/ logic [31:0] value_bits_5;
wire [31:0] _527 = values[4];
/*mux_wire*/ logic [31:0] _525_value;
wire [31:0] _525_bits;
wire  _529 = value_bits_5[0];
wire  _533 = value_bits_5[1];
wire  _537 = value_bits_5[2];
wire  _541 = value_bits_5[3];
wire  _545 = value_bits_5[4];
wire  _549 = value_bits_5[5];
wire  _553 = value_bits_5[6];
wire  _557 = value_bits_5[7];
wire  _561 = value_bits_5[8];
wire  _565 = value_bits_5[9];
wire  _569 = value_bits_5[10];
wire  _573 = value_bits_5[11];
wire  _577 = value_bits_5[12];
wire  _581 = value_bits_5[13];
wire  _585 = value_bits_5[14];
wire  _589 = value_bits_5[15];
wire  _593 = value_bits_5[16];
wire  _597 = value_bits_5[17];
wire  _601 = value_bits_5[18];
wire  _605 = value_bits_5[19];
wire  _609 = value_bits_5[20];
wire  _613 = value_bits_5[21];
wire  _617 = value_bits_5[22];
wire  _621 = value_bits_5[23];
wire  _625 = value_bits_5[24];
wire  _629 = value_bits_5[25];
wire  _633 = value_bits_5[26];
wire  _637 = value_bits_5[27];
wire  _641 = value_bits_5[28];
wire  _645 = value_bits_5[29];
wire  _649 = value_bits_5[30];
wire  _653 = value_bits_5[31];
/*mux_wire*/ logic [31:0] value_bits_6;
wire [31:0] _658 = values[5];
/*mux_wire*/ logic [31:0] _656_value;
wire [31:0] _656_bits;
wire  _660 = value_bits_6[0];
wire  _664 = value_bits_6[1];
wire  _668 = value_bits_6[2];
wire  _672 = value_bits_6[3];
wire  _676 = value_bits_6[4];
wire  _680 = value_bits_6[5];
wire  _684 = value_bits_6[6];
wire  _688 = value_bits_6[7];
wire  _692 = value_bits_6[8];
wire  _696 = value_bits_6[9];
wire  _700 = value_bits_6[10];
wire  _704 = value_bits_6[11];
wire  _708 = value_bits_6[12];
wire  _712 = value_bits_6[13];
wire  _716 = value_bits_6[14];
wire  _720 = value_bits_6[15];
wire  _724 = value_bits_6[16];
wire  _728 = value_bits_6[17];
wire  _732 = value_bits_6[18];
wire  _736 = value_bits_6[19];
wire  _740 = value_bits_6[20];
wire  _744 = value_bits_6[21];
wire  _748 = value_bits_6[22];
wire  _752 = value_bits_6[23];
wire  _756 = value_bits_6[24];
wire  _760 = value_bits_6[25];
wire  _764 = value_bits_6[26];
wire  _768 = value_bits_6[27];
wire  _772 = value_bits_6[28];
wire  _776 = value_bits_6[29];
wire  _780 = value_bits_6[30];
wire  _784 = value_bits_6[31];
/*mux_wire*/ logic [31:0] value_bits_7;
wire [31:0] _789 = values[6];
/*mux_wire*/ logic [31:0] _787_value;
wire [31:0] _787_bits;
wire  _791 = value_bits_7[0];
wire  _795 = value_bits_7[1];
wire  _799 = value_bits_7[2];
wire  _803 = value_bits_7[3];
wire  _807 = value_bits_7[4];
wire  _811 = value_bits_7[5];
wire  _815 = value_bits_7[6];
wire  _819 = value_bits_7[7];
wire  _823 = value_bits_7[8];
wire  _827 = value_bits_7[9];
wire  _831 = value_bits_7[10];
wire  _835 = value_bits_7[11];
wire  _839 = value_bits_7[12];
wire  _843 = value_bits_7[13];
wire  _847 = value_bits_7[14];
wire  _851 = value_bits_7[15];
wire  _855 = value_bits_7[16];
wire  _859 = value_bits_7[17];
wire  _863 = value_bits_7[18];
wire  _867 = value_bits_7[19];
wire  _871 = value_bits_7[20];
wire  _875 = value_bits_7[21];
wire  _879 = value_bits_7[22];
wire  _883 = value_bits_7[23];
wire  _887 = value_bits_7[24];
wire  _891 = value_bits_7[25];
wire  _895 = value_bits_7[26];
wire  _899 = value_bits_7[27];
wire  _903 = value_bits_7[28];
wire  _907 = value_bits_7[29];
wire  _911 = value_bits_7[30];
wire  _915 = value_bits_7[31];
/*mux_wire*/ logic [31:0] value_bits_8;
wire [31:0] _920 = values[7];
/*mux_wire*/ logic [31:0] _918_value;
wire [31:0] _918_bits;
wire  _922 = value_bits_8[0];
wire  _926 = value_bits_8[1];
wire  _930 = value_bits_8[2];
wire  _934 = value_bits_8[3];
wire  _938 = value_bits_8[4];
wire  _942 = value_bits_8[5];
wire  _946 = value_bits_8[6];
wire  _950 = value_bits_8[7];
wire  _954 = value_bits_8[8];
wire  _958 = value_bits_8[9];
wire  _962 = value_bits_8[10];
wire  _966 = value_bits_8[11];
wire  _970 = value_bits_8[12];
wire  _974 = value_bits_8[13];
wire  _978 = value_bits_8[14];
wire  _982 = value_bits_8[15];
wire  _986 = value_bits_8[16];
wire  _990 = value_bits_8[17];
wire  _994 = value_bits_8[18];
wire  _998 = value_bits_8[19];
wire  _1002 = value_bits_8[20];
wire  _1006 = value_bits_8[21];
wire  _1010 = value_bits_8[22];
wire  _1014 = value_bits_8[23];
wire  _1018 = value_bits_8[24];
wire  _1022 = value_bits_8[25];
wire  _1026 = value_bits_8[26];
wire  _1030 = value_bits_8[27];
wire  _1034 = value_bits_8[28];
wire  _1038 = value_bits_8[29];
wire  _1042 = value_bits_8[30];
wire  _1046 = value_bits_8[31];
/*mux_wire*/ logic [31:0] value_bits_9;
wire [31:0] _1051 = values[8];
/*mux_wire*/ logic [31:0] _1049_value;
wire [31:0] _1049_bits;
wire  _1053 = value_bits_9[0];
wire  _1057 = value_bits_9[1];
wire  _1061 = value_bits_9[2];
wire  _1065 = value_bits_9[3];
wire  _1069 = value_bits_9[4];
wire  _1073 = value_bits_9[5];
wire  _1077 = value_bits_9[6];
wire  _1081 = value_bits_9[7];
wire  _1085 = value_bits_9[8];
wire  _1089 = value_bits_9[9];
wire  _1093 = value_bits_9[10];
wire  _1097 = value_bits_9[11];
wire  _1101 = value_bits_9[12];
wire  _1105 = value_bits_9[13];
wire  _1109 = value_bits_9[14];
wire  _1113 = value_bits_9[15];
wire  _1117 = value_bits_9[16];
wire  _1121 = value_bits_9[17];
wire  _1125 = value_bits_9[18];
wire  _1129 = value_bits_9[19];
wire  _1133 = value_bits_9[20];
wire  _1137 = value_bits_9[21];
wire  _1141 = value_bits_9[22];
wire  _1145 = value_bits_9[23];
wire  _1149 = value_bits_9[24];
wire  _1153 = value_bits_9[25];
wire  _1157 = value_bits_9[26];
wire  _1161 = value_bits_9[27];
wire  _1165 = value_bits_9[28];
wire  _1169 = value_bits_9[29];
wire  _1173 = value_bits_9[30];
wire  _1177 = value_bits_9[31];
/*mux_wire*/ logic [31:0] value_bits_10;
wire [31:0] _1182 = values[9];
/*mux_wire*/ logic [31:0] _1180_value;
wire [31:0] _1180_bits;
wire  _1184 = value_bits_10[0];
wire  _1188 = value_bits_10[1];
wire  _1192 = value_bits_10[2];
wire  _1196 = value_bits_10[3];
wire  _1200 = value_bits_10[4];
wire  _1204 = value_bits_10[5];
wire  _1208 = value_bits_10[6];
wire  _1212 = value_bits_10[7];
wire  _1216 = value_bits_10[8];
wire  _1220 = value_bits_10[9];
wire  _1224 = value_bits_10[10];
wire  _1228 = value_bits_10[11];
wire  _1232 = value_bits_10[12];
wire  _1236 = value_bits_10[13];
wire  _1240 = value_bits_10[14];
wire  _1244 = value_bits_10[15];
wire  _1248 = value_bits_10[16];
wire  _1252 = value_bits_10[17];
wire  _1256 = value_bits_10[18];
wire  _1260 = value_bits_10[19];
wire  _1264 = value_bits_10[20];
wire  _1268 = value_bits_10[21];
wire  _1272 = value_bits_10[22];
wire  _1276 = value_bits_10[23];
wire  _1280 = value_bits_10[24];
wire  _1284 = value_bits_10[25];
wire  _1288 = value_bits_10[26];
wire  _1292 = value_bits_10[27];
wire  _1296 = value_bits_10[28];
wire  _1300 = value_bits_10[29];
wire  _1304 = value_bits_10[30];
wire  _1308 = value_bits_10[31];
wire [9:0] _1312 = split_into_bits[0];
wire [9:0] _1315 = split_into_bits[1];
wire [9:0] _1318 = split_into_bits[2];
wire [9:0] _1321 = split_into_bits[3];
wire [9:0] _1324 = split_into_bits[4];
wire [9:0] _1327 = split_into_bits[5];
wire [9:0] _1330 = split_into_bits[6];
wire [9:0] _1333 = split_into_bits[7];
wire [9:0] _1336 = split_into_bits[8];
wire [9:0] _1339 = split_into_bits[9];
wire [9:0] _1342 = split_into_bits[10];
wire [9:0] _1345 = split_into_bits[11];
wire [9:0] _1348 = split_into_bits[12];
wire [9:0] _1351 = split_into_bits[13];
wire [9:0] _1354 = split_into_bits[14];
wire [9:0] _1357 = split_into_bits[15];
wire [9:0] _1360 = split_into_bits[16];
wire [9:0] _1363 = split_into_bits[17];
wire [9:0] _1366 = split_into_bits[18];
wire [9:0] _1369 = split_into_bits[19];
wire [9:0] _1372 = split_into_bits[20];
wire [9:0] _1375 = split_into_bits[21];
wire [9:0] _1378 = split_into_bits[22];
wire [9:0] _1381 = split_into_bits[23];
wire [9:0] _1384 = split_into_bits[24];
wire [9:0] _1387 = split_into_bits[25];
wire [9:0] _1390 = split_into_bits[26];
wire [9:0] _1393 = split_into_bits[27];
wire [9:0] _1396 = split_into_bits[28];
wire [9:0] _1399 = split_into_bits[29];
wire [9:0] _1402 = split_into_bits[30];
wire [9:0] _1405 = split_into_bits[31];
IntToBits _1(
	.clk(clk),
	.value(_1_value),
	.bits(_1_bits)
);
IntToBits _132(
	.clk(clk),
	.value(_132_value),
	.bits(_132_bits)
);
IntToBits _263(
	.clk(clk),
	.value(_263_value),
	.bits(_263_bits)
);
IntToBits _394(
	.clk(clk),
	.value(_394_value),
	.bits(_394_bits)
);
IntToBits _525(
	.clk(clk),
	.value(_525_value),
	.bits(_525_bits)
);
IntToBits _656(
	.clk(clk),
	.value(_656_value),
	.bits(_656_bits)
);
IntToBits _787(
	.clk(clk),
	.value(_787_value),
	.bits(_787_bits)
);
IntToBits _918(
	.clk(clk),
	.value(_918_value),
	.bits(_918_bits)
);
IntToBits _1049(
	.clk(clk),
	.value(_1049_value),
	.bits(_1049_bits)
);
IntToBits _1180(
	.clk(clk),
	.value(_1180_value),
	.bits(_1180_bits)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	bits[0] = 'x;
	bits[1] = 'x;
	bits[2] = 'x;
	bits[3] = 'x;
	bits[4] = 'x;
	bits[5] = 'x;
	bits[6] = 'x;
	bits[7] = 'x;
	bits[8] = 'x;
	bits[9] = 'x;
	if(shift) bits = _1405;
end
always_ff @(posedge clk) begin
	if(start) split_into_bits[0][0] <= _5;
	if(start) split_into_bits[1][0] <= _9;
	if(start) split_into_bits[2][0] <= _13;
	if(start) split_into_bits[3][0] <= _17;
	if(start) split_into_bits[4][0] <= _21;
	if(start) split_into_bits[5][0] <= _25;
	if(start) split_into_bits[6][0] <= _29;
	if(start) split_into_bits[7][0] <= _33;
	if(start) split_into_bits[8][0] <= _37;
	if(start) split_into_bits[9][0] <= _41;
	if(start) split_into_bits[10][0] <= _45;
	if(start) split_into_bits[11][0] <= _49;
	if(start) split_into_bits[12][0] <= _53;
	if(start) split_into_bits[13][0] <= _57;
	if(start) split_into_bits[14][0] <= _61;
	if(start) split_into_bits[15][0] <= _65;
	if(start) split_into_bits[16][0] <= _69;
	if(start) split_into_bits[17][0] <= _73;
	if(start) split_into_bits[18][0] <= _77;
	if(start) split_into_bits[19][0] <= _81;
	if(start) split_into_bits[20][0] <= _85;
	if(start) split_into_bits[21][0] <= _89;
	if(start) split_into_bits[22][0] <= _93;
	if(start) split_into_bits[23][0] <= _97;
	if(start) split_into_bits[24][0] <= _101;
	if(start) split_into_bits[25][0] <= _105;
	if(start) split_into_bits[26][0] <= _109;
	if(start) split_into_bits[27][0] <= _113;
	if(start) split_into_bits[28][0] <= _117;
	if(start) split_into_bits[29][0] <= _121;
	if(start) split_into_bits[30][0] <= _125;
	if(start) split_into_bits[31][0] <= _129;
	if(start) split_into_bits[0][1] <= _136;
	if(start) split_into_bits[1][1] <= _140;
	if(start) split_into_bits[2][1] <= _144;
	if(start) split_into_bits[3][1] <= _148;
	if(start) split_into_bits[4][1] <= _152;
	if(start) split_into_bits[5][1] <= _156;
	if(start) split_into_bits[6][1] <= _160;
	if(start) split_into_bits[7][1] <= _164;
	if(start) split_into_bits[8][1] <= _168;
	if(start) split_into_bits[9][1] <= _172;
	if(start) split_into_bits[10][1] <= _176;
	if(start) split_into_bits[11][1] <= _180;
	if(start) split_into_bits[12][1] <= _184;
	if(start) split_into_bits[13][1] <= _188;
	if(start) split_into_bits[14][1] <= _192;
	if(start) split_into_bits[15][1] <= _196;
	if(start) split_into_bits[16][1] <= _200;
	if(start) split_into_bits[17][1] <= _204;
	if(start) split_into_bits[18][1] <= _208;
	if(start) split_into_bits[19][1] <= _212;
	if(start) split_into_bits[20][1] <= _216;
	if(start) split_into_bits[21][1] <= _220;
	if(start) split_into_bits[22][1] <= _224;
	if(start) split_into_bits[23][1] <= _228;
	if(start) split_into_bits[24][1] <= _232;
	if(start) split_into_bits[25][1] <= _236;
	if(start) split_into_bits[26][1] <= _240;
	if(start) split_into_bits[27][1] <= _244;
	if(start) split_into_bits[28][1] <= _248;
	if(start) split_into_bits[29][1] <= _252;
	if(start) split_into_bits[30][1] <= _256;
	if(start) split_into_bits[31][1] <= _260;
	if(start) split_into_bits[0][2] <= _267;
	if(start) split_into_bits[1][2] <= _271;
	if(start) split_into_bits[2][2] <= _275;
	if(start) split_into_bits[3][2] <= _279;
	if(start) split_into_bits[4][2] <= _283;
	if(start) split_into_bits[5][2] <= _287;
	if(start) split_into_bits[6][2] <= _291;
	if(start) split_into_bits[7][2] <= _295;
	if(start) split_into_bits[8][2] <= _299;
	if(start) split_into_bits[9][2] <= _303;
	if(start) split_into_bits[10][2] <= _307;
	if(start) split_into_bits[11][2] <= _311;
	if(start) split_into_bits[12][2] <= _315;
	if(start) split_into_bits[13][2] <= _319;
	if(start) split_into_bits[14][2] <= _323;
	if(start) split_into_bits[15][2] <= _327;
	if(start) split_into_bits[16][2] <= _331;
	if(start) split_into_bits[17][2] <= _335;
	if(start) split_into_bits[18][2] <= _339;
	if(start) split_into_bits[19][2] <= _343;
	if(start) split_into_bits[20][2] <= _347;
	if(start) split_into_bits[21][2] <= _351;
	if(start) split_into_bits[22][2] <= _355;
	if(start) split_into_bits[23][2] <= _359;
	if(start) split_into_bits[24][2] <= _363;
	if(start) split_into_bits[25][2] <= _367;
	if(start) split_into_bits[26][2] <= _371;
	if(start) split_into_bits[27][2] <= _375;
	if(start) split_into_bits[28][2] <= _379;
	if(start) split_into_bits[29][2] <= _383;
	if(start) split_into_bits[30][2] <= _387;
	if(start) split_into_bits[31][2] <= _391;
	if(start) split_into_bits[0][3] <= _398;
	if(start) split_into_bits[1][3] <= _402;
	if(start) split_into_bits[2][3] <= _406;
	if(start) split_into_bits[3][3] <= _410;
	if(start) split_into_bits[4][3] <= _414;
	if(start) split_into_bits[5][3] <= _418;
	if(start) split_into_bits[6][3] <= _422;
	if(start) split_into_bits[7][3] <= _426;
	if(start) split_into_bits[8][3] <= _430;
	if(start) split_into_bits[9][3] <= _434;
	if(start) split_into_bits[10][3] <= _438;
	if(start) split_into_bits[11][3] <= _442;
	if(start) split_into_bits[12][3] <= _446;
	if(start) split_into_bits[13][3] <= _450;
	if(start) split_into_bits[14][3] <= _454;
	if(start) split_into_bits[15][3] <= _458;
	if(start) split_into_bits[16][3] <= _462;
	if(start) split_into_bits[17][3] <= _466;
	if(start) split_into_bits[18][3] <= _470;
	if(start) split_into_bits[19][3] <= _474;
	if(start) split_into_bits[20][3] <= _478;
	if(start) split_into_bits[21][3] <= _482;
	if(start) split_into_bits[22][3] <= _486;
	if(start) split_into_bits[23][3] <= _490;
	if(start) split_into_bits[24][3] <= _494;
	if(start) split_into_bits[25][3] <= _498;
	if(start) split_into_bits[26][3] <= _502;
	if(start) split_into_bits[27][3] <= _506;
	if(start) split_into_bits[28][3] <= _510;
	if(start) split_into_bits[29][3] <= _514;
	if(start) split_into_bits[30][3] <= _518;
	if(start) split_into_bits[31][3] <= _522;
	if(start) split_into_bits[0][4] <= _529;
	if(start) split_into_bits[1][4] <= _533;
	if(start) split_into_bits[2][4] <= _537;
	if(start) split_into_bits[3][4] <= _541;
	if(start) split_into_bits[4][4] <= _545;
	if(start) split_into_bits[5][4] <= _549;
	if(start) split_into_bits[6][4] <= _553;
	if(start) split_into_bits[7][4] <= _557;
	if(start) split_into_bits[8][4] <= _561;
	if(start) split_into_bits[9][4] <= _565;
	if(start) split_into_bits[10][4] <= _569;
	if(start) split_into_bits[11][4] <= _573;
	if(start) split_into_bits[12][4] <= _577;
	if(start) split_into_bits[13][4] <= _581;
	if(start) split_into_bits[14][4] <= _585;
	if(start) split_into_bits[15][4] <= _589;
	if(start) split_into_bits[16][4] <= _593;
	if(start) split_into_bits[17][4] <= _597;
	if(start) split_into_bits[18][4] <= _601;
	if(start) split_into_bits[19][4] <= _605;
	if(start) split_into_bits[20][4] <= _609;
	if(start) split_into_bits[21][4] <= _613;
	if(start) split_into_bits[22][4] <= _617;
	if(start) split_into_bits[23][4] <= _621;
	if(start) split_into_bits[24][4] <= _625;
	if(start) split_into_bits[25][4] <= _629;
	if(start) split_into_bits[26][4] <= _633;
	if(start) split_into_bits[27][4] <= _637;
	if(start) split_into_bits[28][4] <= _641;
	if(start) split_into_bits[29][4] <= _645;
	if(start) split_into_bits[30][4] <= _649;
	if(start) split_into_bits[31][4] <= _653;
	if(start) split_into_bits[0][5] <= _660;
	if(start) split_into_bits[1][5] <= _664;
	if(start) split_into_bits[2][5] <= _668;
	if(start) split_into_bits[3][5] <= _672;
	if(start) split_into_bits[4][5] <= _676;
	if(start) split_into_bits[5][5] <= _680;
	if(start) split_into_bits[6][5] <= _684;
	if(start) split_into_bits[7][5] <= _688;
	if(start) split_into_bits[8][5] <= _692;
	if(start) split_into_bits[9][5] <= _696;
	if(start) split_into_bits[10][5] <= _700;
	if(start) split_into_bits[11][5] <= _704;
	if(start) split_into_bits[12][5] <= _708;
	if(start) split_into_bits[13][5] <= _712;
	if(start) split_into_bits[14][5] <= _716;
	if(start) split_into_bits[15][5] <= _720;
	if(start) split_into_bits[16][5] <= _724;
	if(start) split_into_bits[17][5] <= _728;
	if(start) split_into_bits[18][5] <= _732;
	if(start) split_into_bits[19][5] <= _736;
	if(start) split_into_bits[20][5] <= _740;
	if(start) split_into_bits[21][5] <= _744;
	if(start) split_into_bits[22][5] <= _748;
	if(start) split_into_bits[23][5] <= _752;
	if(start) split_into_bits[24][5] <= _756;
	if(start) split_into_bits[25][5] <= _760;
	if(start) split_into_bits[26][5] <= _764;
	if(start) split_into_bits[27][5] <= _768;
	if(start) split_into_bits[28][5] <= _772;
	if(start) split_into_bits[29][5] <= _776;
	if(start) split_into_bits[30][5] <= _780;
	if(start) split_into_bits[31][5] <= _784;
	if(start) split_into_bits[0][6] <= _791;
	if(start) split_into_bits[1][6] <= _795;
	if(start) split_into_bits[2][6] <= _799;
	if(start) split_into_bits[3][6] <= _803;
	if(start) split_into_bits[4][6] <= _807;
	if(start) split_into_bits[5][6] <= _811;
	if(start) split_into_bits[6][6] <= _815;
	if(start) split_into_bits[7][6] <= _819;
	if(start) split_into_bits[8][6] <= _823;
	if(start) split_into_bits[9][6] <= _827;
	if(start) split_into_bits[10][6] <= _831;
	if(start) split_into_bits[11][6] <= _835;
	if(start) split_into_bits[12][6] <= _839;
	if(start) split_into_bits[13][6] <= _843;
	if(start) split_into_bits[14][6] <= _847;
	if(start) split_into_bits[15][6] <= _851;
	if(start) split_into_bits[16][6] <= _855;
	if(start) split_into_bits[17][6] <= _859;
	if(start) split_into_bits[18][6] <= _863;
	if(start) split_into_bits[19][6] <= _867;
	if(start) split_into_bits[20][6] <= _871;
	if(start) split_into_bits[21][6] <= _875;
	if(start) split_into_bits[22][6] <= _879;
	if(start) split_into_bits[23][6] <= _883;
	if(start) split_into_bits[24][6] <= _887;
	if(start) split_into_bits[25][6] <= _891;
	if(start) split_into_bits[26][6] <= _895;
	if(start) split_into_bits[27][6] <= _899;
	if(start) split_into_bits[28][6] <= _903;
	if(start) split_into_bits[29][6] <= _907;
	if(start) split_into_bits[30][6] <= _911;
	if(start) split_into_bits[31][6] <= _915;
	if(start) split_into_bits[0][7] <= _922;
	if(start) split_into_bits[1][7] <= _926;
	if(start) split_into_bits[2][7] <= _930;
	if(start) split_into_bits[3][7] <= _934;
	if(start) split_into_bits[4][7] <= _938;
	if(start) split_into_bits[5][7] <= _942;
	if(start) split_into_bits[6][7] <= _946;
	if(start) split_into_bits[7][7] <= _950;
	if(start) split_into_bits[8][7] <= _954;
	if(start) split_into_bits[9][7] <= _958;
	if(start) split_into_bits[10][7] <= _962;
	if(start) split_into_bits[11][7] <= _966;
	if(start) split_into_bits[12][7] <= _970;
	if(start) split_into_bits[13][7] <= _974;
	if(start) split_into_bits[14][7] <= _978;
	if(start) split_into_bits[15][7] <= _982;
	if(start) split_into_bits[16][7] <= _986;
	if(start) split_into_bits[17][7] <= _990;
	if(start) split_into_bits[18][7] <= _994;
	if(start) split_into_bits[19][7] <= _998;
	if(start) split_into_bits[20][7] <= _1002;
	if(start) split_into_bits[21][7] <= _1006;
	if(start) split_into_bits[22][7] <= _1010;
	if(start) split_into_bits[23][7] <= _1014;
	if(start) split_into_bits[24][7] <= _1018;
	if(start) split_into_bits[25][7] <= _1022;
	if(start) split_into_bits[26][7] <= _1026;
	if(start) split_into_bits[27][7] <= _1030;
	if(start) split_into_bits[28][7] <= _1034;
	if(start) split_into_bits[29][7] <= _1038;
	if(start) split_into_bits[30][7] <= _1042;
	if(start) split_into_bits[31][7] <= _1046;
	if(start) split_into_bits[0][8] <= _1053;
	if(start) split_into_bits[1][8] <= _1057;
	if(start) split_into_bits[2][8] <= _1061;
	if(start) split_into_bits[3][8] <= _1065;
	if(start) split_into_bits[4][8] <= _1069;
	if(start) split_into_bits[5][8] <= _1073;
	if(start) split_into_bits[6][8] <= _1077;
	if(start) split_into_bits[7][8] <= _1081;
	if(start) split_into_bits[8][8] <= _1085;
	if(start) split_into_bits[9][8] <= _1089;
	if(start) split_into_bits[10][8] <= _1093;
	if(start) split_into_bits[11][8] <= _1097;
	if(start) split_into_bits[12][8] <= _1101;
	if(start) split_into_bits[13][8] <= _1105;
	if(start) split_into_bits[14][8] <= _1109;
	if(start) split_into_bits[15][8] <= _1113;
	if(start) split_into_bits[16][8] <= _1117;
	if(start) split_into_bits[17][8] <= _1121;
	if(start) split_into_bits[18][8] <= _1125;
	if(start) split_into_bits[19][8] <= _1129;
	if(start) split_into_bits[20][8] <= _1133;
	if(start) split_into_bits[21][8] <= _1137;
	if(start) split_into_bits[22][8] <= _1141;
	if(start) split_into_bits[23][8] <= _1145;
	if(start) split_into_bits[24][8] <= _1149;
	if(start) split_into_bits[25][8] <= _1153;
	if(start) split_into_bits[26][8] <= _1157;
	if(start) split_into_bits[27][8] <= _1161;
	if(start) split_into_bits[28][8] <= _1165;
	if(start) split_into_bits[29][8] <= _1169;
	if(start) split_into_bits[30][8] <= _1173;
	if(start) split_into_bits[31][8] <= _1177;
	if(start) split_into_bits[0][9] <= _1184;
	if(start) split_into_bits[1][9] <= _1188;
	if(start) split_into_bits[2][9] <= _1192;
	if(start) split_into_bits[3][9] <= _1196;
	if(start) split_into_bits[4][9] <= _1200;
	if(start) split_into_bits[5][9] <= _1204;
	if(start) split_into_bits[6][9] <= _1208;
	if(start) split_into_bits[7][9] <= _1212;
	if(start) split_into_bits[8][9] <= _1216;
	if(start) split_into_bits[9][9] <= _1220;
	if(start) split_into_bits[10][9] <= _1224;
	if(start) split_into_bits[11][9] <= _1228;
	if(start) split_into_bits[12][9] <= _1232;
	if(start) split_into_bits[13][9] <= _1236;
	if(start) split_into_bits[14][9] <= _1240;
	if(start) split_into_bits[15][9] <= _1244;
	if(start) split_into_bits[16][9] <= _1248;
	if(start) split_into_bits[17][9] <= _1252;
	if(start) split_into_bits[18][9] <= _1256;
	if(start) split_into_bits[19][9] <= _1260;
	if(start) split_into_bits[20][9] <= _1264;
	if(start) split_into_bits[21][9] <= _1268;
	if(start) split_into_bits[22][9] <= _1272;
	if(start) split_into_bits[23][9] <= _1276;
	if(start) split_into_bits[24][9] <= _1280;
	if(start) split_into_bits[25][9] <= _1284;
	if(start) split_into_bits[26][9] <= _1288;
	if(start) split_into_bits[27][9] <= _1292;
	if(start) split_into_bits[28][9] <= _1296;
	if(start) split_into_bits[29][9] <= _1300;
	if(start) split_into_bits[30][9] <= _1304;
	if(start) split_into_bits[31][9] <= _1308;
	if(!start) if(shift) split_into_bits[1] <= _1312;
	if(!start) if(shift) split_into_bits[2] <= _1315;
	if(!start) if(shift) split_into_bits[3] <= _1318;
	if(!start) if(shift) split_into_bits[4] <= _1321;
	if(!start) if(shift) split_into_bits[5] <= _1324;
	if(!start) if(shift) split_into_bits[6] <= _1327;
	if(!start) if(shift) split_into_bits[7] <= _1330;
	if(!start) if(shift) split_into_bits[8] <= _1333;
	if(!start) if(shift) split_into_bits[9] <= _1336;
	if(!start) if(shift) split_into_bits[10] <= _1339;
	if(!start) if(shift) split_into_bits[11] <= _1342;
	if(!start) if(shift) split_into_bits[12] <= _1345;
	if(!start) if(shift) split_into_bits[13] <= _1348;
	if(!start) if(shift) split_into_bits[14] <= _1351;
	if(!start) if(shift) split_into_bits[15] <= _1354;
	if(!start) if(shift) split_into_bits[16] <= _1357;
	if(!start) if(shift) split_into_bits[17] <= _1360;
	if(!start) if(shift) split_into_bits[18] <= _1363;
	if(!start) if(shift) split_into_bits[19] <= _1366;
	if(!start) if(shift) split_into_bits[20] <= _1369;
	if(!start) if(shift) split_into_bits[21] <= _1372;
	if(!start) if(shift) split_into_bits[22] <= _1375;
	if(!start) if(shift) split_into_bits[23] <= _1378;
	if(!start) if(shift) split_into_bits[24] <= _1381;
	if(!start) if(shift) split_into_bits[25] <= _1384;
	if(!start) if(shift) split_into_bits[26] <= _1387;
	if(!start) if(shift) split_into_bits[27] <= _1390;
	if(!start) if(shift) split_into_bits[28] <= _1393;
	if(!start) if(shift) split_into_bits[29] <= _1396;
	if(!start) if(shift) split_into_bits[30] <= _1399;
	if(!start) if(shift) split_into_bits[31] <= _1402;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits[0] = 'x;
	value_bits[1] = 'x;
	value_bits[2] = 'x;
	value_bits[3] = 'x;
	value_bits[4] = 'x;
	value_bits[5] = 'x;
	value_bits[6] = 'x;
	value_bits[7] = 'x;
	value_bits[8] = 'x;
	value_bits[9] = 'x;
	value_bits[10] = 'x;
	value_bits[11] = 'x;
	value_bits[12] = 'x;
	value_bits[13] = 'x;
	value_bits[14] = 'x;
	value_bits[15] = 'x;
	value_bits[16] = 'x;
	value_bits[17] = 'x;
	value_bits[18] = 'x;
	value_bits[19] = 'x;
	value_bits[20] = 'x;
	value_bits[21] = 'x;
	value_bits[22] = 'x;
	value_bits[23] = 'x;
	value_bits[24] = 'x;
	value_bits[25] = 'x;
	value_bits[26] = 'x;
	value_bits[27] = 'x;
	value_bits[28] = 'x;
	value_bits[29] = 'x;
	value_bits[30] = 'x;
	value_bits[31] = 'x;
	if(start) value_bits = _1_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1_value = 'x;
	if(start) _1_value = _3;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_2[0] = 'x;
	value_bits_2[1] = 'x;
	value_bits_2[2] = 'x;
	value_bits_2[3] = 'x;
	value_bits_2[4] = 'x;
	value_bits_2[5] = 'x;
	value_bits_2[6] = 'x;
	value_bits_2[7] = 'x;
	value_bits_2[8] = 'x;
	value_bits_2[9] = 'x;
	value_bits_2[10] = 'x;
	value_bits_2[11] = 'x;
	value_bits_2[12] = 'x;
	value_bits_2[13] = 'x;
	value_bits_2[14] = 'x;
	value_bits_2[15] = 'x;
	value_bits_2[16] = 'x;
	value_bits_2[17] = 'x;
	value_bits_2[18] = 'x;
	value_bits_2[19] = 'x;
	value_bits_2[20] = 'x;
	value_bits_2[21] = 'x;
	value_bits_2[22] = 'x;
	value_bits_2[23] = 'x;
	value_bits_2[24] = 'x;
	value_bits_2[25] = 'x;
	value_bits_2[26] = 'x;
	value_bits_2[27] = 'x;
	value_bits_2[28] = 'x;
	value_bits_2[29] = 'x;
	value_bits_2[30] = 'x;
	value_bits_2[31] = 'x;
	if(start) value_bits_2 = _132_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_132_value = 'x;
	if(start) _132_value = _134;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_3[0] = 'x;
	value_bits_3[1] = 'x;
	value_bits_3[2] = 'x;
	value_bits_3[3] = 'x;
	value_bits_3[4] = 'x;
	value_bits_3[5] = 'x;
	value_bits_3[6] = 'x;
	value_bits_3[7] = 'x;
	value_bits_3[8] = 'x;
	value_bits_3[9] = 'x;
	value_bits_3[10] = 'x;
	value_bits_3[11] = 'x;
	value_bits_3[12] = 'x;
	value_bits_3[13] = 'x;
	value_bits_3[14] = 'x;
	value_bits_3[15] = 'x;
	value_bits_3[16] = 'x;
	value_bits_3[17] = 'x;
	value_bits_3[18] = 'x;
	value_bits_3[19] = 'x;
	value_bits_3[20] = 'x;
	value_bits_3[21] = 'x;
	value_bits_3[22] = 'x;
	value_bits_3[23] = 'x;
	value_bits_3[24] = 'x;
	value_bits_3[25] = 'x;
	value_bits_3[26] = 'x;
	value_bits_3[27] = 'x;
	value_bits_3[28] = 'x;
	value_bits_3[29] = 'x;
	value_bits_3[30] = 'x;
	value_bits_3[31] = 'x;
	if(start) value_bits_3 = _263_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_263_value = 'x;
	if(start) _263_value = _265;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_4[0] = 'x;
	value_bits_4[1] = 'x;
	value_bits_4[2] = 'x;
	value_bits_4[3] = 'x;
	value_bits_4[4] = 'x;
	value_bits_4[5] = 'x;
	value_bits_4[6] = 'x;
	value_bits_4[7] = 'x;
	value_bits_4[8] = 'x;
	value_bits_4[9] = 'x;
	value_bits_4[10] = 'x;
	value_bits_4[11] = 'x;
	value_bits_4[12] = 'x;
	value_bits_4[13] = 'x;
	value_bits_4[14] = 'x;
	value_bits_4[15] = 'x;
	value_bits_4[16] = 'x;
	value_bits_4[17] = 'x;
	value_bits_4[18] = 'x;
	value_bits_4[19] = 'x;
	value_bits_4[20] = 'x;
	value_bits_4[21] = 'x;
	value_bits_4[22] = 'x;
	value_bits_4[23] = 'x;
	value_bits_4[24] = 'x;
	value_bits_4[25] = 'x;
	value_bits_4[26] = 'x;
	value_bits_4[27] = 'x;
	value_bits_4[28] = 'x;
	value_bits_4[29] = 'x;
	value_bits_4[30] = 'x;
	value_bits_4[31] = 'x;
	if(start) value_bits_4 = _394_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_394_value = 'x;
	if(start) _394_value = _396;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_5[0] = 'x;
	value_bits_5[1] = 'x;
	value_bits_5[2] = 'x;
	value_bits_5[3] = 'x;
	value_bits_5[4] = 'x;
	value_bits_5[5] = 'x;
	value_bits_5[6] = 'x;
	value_bits_5[7] = 'x;
	value_bits_5[8] = 'x;
	value_bits_5[9] = 'x;
	value_bits_5[10] = 'x;
	value_bits_5[11] = 'x;
	value_bits_5[12] = 'x;
	value_bits_5[13] = 'x;
	value_bits_5[14] = 'x;
	value_bits_5[15] = 'x;
	value_bits_5[16] = 'x;
	value_bits_5[17] = 'x;
	value_bits_5[18] = 'x;
	value_bits_5[19] = 'x;
	value_bits_5[20] = 'x;
	value_bits_5[21] = 'x;
	value_bits_5[22] = 'x;
	value_bits_5[23] = 'x;
	value_bits_5[24] = 'x;
	value_bits_5[25] = 'x;
	value_bits_5[26] = 'x;
	value_bits_5[27] = 'x;
	value_bits_5[28] = 'x;
	value_bits_5[29] = 'x;
	value_bits_5[30] = 'x;
	value_bits_5[31] = 'x;
	if(start) value_bits_5 = _525_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_525_value = 'x;
	if(start) _525_value = _527;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_6[0] = 'x;
	value_bits_6[1] = 'x;
	value_bits_6[2] = 'x;
	value_bits_6[3] = 'x;
	value_bits_6[4] = 'x;
	value_bits_6[5] = 'x;
	value_bits_6[6] = 'x;
	value_bits_6[7] = 'x;
	value_bits_6[8] = 'x;
	value_bits_6[9] = 'x;
	value_bits_6[10] = 'x;
	value_bits_6[11] = 'x;
	value_bits_6[12] = 'x;
	value_bits_6[13] = 'x;
	value_bits_6[14] = 'x;
	value_bits_6[15] = 'x;
	value_bits_6[16] = 'x;
	value_bits_6[17] = 'x;
	value_bits_6[18] = 'x;
	value_bits_6[19] = 'x;
	value_bits_6[20] = 'x;
	value_bits_6[21] = 'x;
	value_bits_6[22] = 'x;
	value_bits_6[23] = 'x;
	value_bits_6[24] = 'x;
	value_bits_6[25] = 'x;
	value_bits_6[26] = 'x;
	value_bits_6[27] = 'x;
	value_bits_6[28] = 'x;
	value_bits_6[29] = 'x;
	value_bits_6[30] = 'x;
	value_bits_6[31] = 'x;
	if(start) value_bits_6 = _656_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_656_value = 'x;
	if(start) _656_value = _658;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_7[0] = 'x;
	value_bits_7[1] = 'x;
	value_bits_7[2] = 'x;
	value_bits_7[3] = 'x;
	value_bits_7[4] = 'x;
	value_bits_7[5] = 'x;
	value_bits_7[6] = 'x;
	value_bits_7[7] = 'x;
	value_bits_7[8] = 'x;
	value_bits_7[9] = 'x;
	value_bits_7[10] = 'x;
	value_bits_7[11] = 'x;
	value_bits_7[12] = 'x;
	value_bits_7[13] = 'x;
	value_bits_7[14] = 'x;
	value_bits_7[15] = 'x;
	value_bits_7[16] = 'x;
	value_bits_7[17] = 'x;
	value_bits_7[18] = 'x;
	value_bits_7[19] = 'x;
	value_bits_7[20] = 'x;
	value_bits_7[21] = 'x;
	value_bits_7[22] = 'x;
	value_bits_7[23] = 'x;
	value_bits_7[24] = 'x;
	value_bits_7[25] = 'x;
	value_bits_7[26] = 'x;
	value_bits_7[27] = 'x;
	value_bits_7[28] = 'x;
	value_bits_7[29] = 'x;
	value_bits_7[30] = 'x;
	value_bits_7[31] = 'x;
	if(start) value_bits_7 = _787_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_787_value = 'x;
	if(start) _787_value = _789;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_8[0] = 'x;
	value_bits_8[1] = 'x;
	value_bits_8[2] = 'x;
	value_bits_8[3] = 'x;
	value_bits_8[4] = 'x;
	value_bits_8[5] = 'x;
	value_bits_8[6] = 'x;
	value_bits_8[7] = 'x;
	value_bits_8[8] = 'x;
	value_bits_8[9] = 'x;
	value_bits_8[10] = 'x;
	value_bits_8[11] = 'x;
	value_bits_8[12] = 'x;
	value_bits_8[13] = 'x;
	value_bits_8[14] = 'x;
	value_bits_8[15] = 'x;
	value_bits_8[16] = 'x;
	value_bits_8[17] = 'x;
	value_bits_8[18] = 'x;
	value_bits_8[19] = 'x;
	value_bits_8[20] = 'x;
	value_bits_8[21] = 'x;
	value_bits_8[22] = 'x;
	value_bits_8[23] = 'x;
	value_bits_8[24] = 'x;
	value_bits_8[25] = 'x;
	value_bits_8[26] = 'x;
	value_bits_8[27] = 'x;
	value_bits_8[28] = 'x;
	value_bits_8[29] = 'x;
	value_bits_8[30] = 'x;
	value_bits_8[31] = 'x;
	if(start) value_bits_8 = _918_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_918_value = 'x;
	if(start) _918_value = _920;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_9[0] = 'x;
	value_bits_9[1] = 'x;
	value_bits_9[2] = 'x;
	value_bits_9[3] = 'x;
	value_bits_9[4] = 'x;
	value_bits_9[5] = 'x;
	value_bits_9[6] = 'x;
	value_bits_9[7] = 'x;
	value_bits_9[8] = 'x;
	value_bits_9[9] = 'x;
	value_bits_9[10] = 'x;
	value_bits_9[11] = 'x;
	value_bits_9[12] = 'x;
	value_bits_9[13] = 'x;
	value_bits_9[14] = 'x;
	value_bits_9[15] = 'x;
	value_bits_9[16] = 'x;
	value_bits_9[17] = 'x;
	value_bits_9[18] = 'x;
	value_bits_9[19] = 'x;
	value_bits_9[20] = 'x;
	value_bits_9[21] = 'x;
	value_bits_9[22] = 'x;
	value_bits_9[23] = 'x;
	value_bits_9[24] = 'x;
	value_bits_9[25] = 'x;
	value_bits_9[26] = 'x;
	value_bits_9[27] = 'x;
	value_bits_9[28] = 'x;
	value_bits_9[29] = 'x;
	value_bits_9[30] = 'x;
	value_bits_9[31] = 'x;
	if(start) value_bits_9 = _1049_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1049_value = 'x;
	if(start) _1049_value = _1051;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	value_bits_10[0] = 'x;
	value_bits_10[1] = 'x;
	value_bits_10[2] = 'x;
	value_bits_10[3] = 'x;
	value_bits_10[4] = 'x;
	value_bits_10[5] = 'x;
	value_bits_10[6] = 'x;
	value_bits_10[7] = 'x;
	value_bits_10[8] = 'x;
	value_bits_10[9] = 'x;
	value_bits_10[10] = 'x;
	value_bits_10[11] = 'x;
	value_bits_10[12] = 'x;
	value_bits_10[13] = 'x;
	value_bits_10[14] = 'x;
	value_bits_10[15] = 'x;
	value_bits_10[16] = 'x;
	value_bits_10[17] = 'x;
	value_bits_10[18] = 'x;
	value_bits_10[19] = 'x;
	value_bits_10[20] = 'x;
	value_bits_10[21] = 'x;
	value_bits_10[22] = 'x;
	value_bits_10[23] = 'x;
	value_bits_10[24] = 'x;
	value_bits_10[25] = 'x;
	value_bits_10[26] = 'x;
	value_bits_10[27] = 'x;
	value_bits_10[28] = 'x;
	value_bits_10[29] = 'x;
	value_bits_10[30] = 'x;
	value_bits_10[31] = 'x;
	if(start) value_bits_10 = _1180_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1180_value = 'x;
	if(start) _1180_value = _1182;
end
endmodule

// ::BitSerialMatrixMultiplyState::<WIDTH = 10, HEIGHT = 15, MATRIX = [[0, 2, 0, 0, 0, 10, 0, 0, 0, 18], [0, 3, 0, 0, 0, 0, 0, 0, 0, 19], [2, 4, 0, 0, 10, 0, 14, 0, 0, 20], [0, 5, 7, 9, 0, 0, 15, 0, 0, 21], [0, 6, 0, 0, 0, 0, 0, 0, 0, 22], [0, 7, 0, 0, 0, 15, 0, 0, 0, 23], [6, 8, 0, 12, 14, 16, 0, 0, 0, 24], [0, 9, 0, 0, 0, 0, 0, 21, 0, 25], [0, 10, 12, 0, 0, 0, 0, 22, 0, 26], [0, 11, 0, 0, 0, 0, 0, 23, 0, 27], [10, 12, 14, 0, 18, 0, 0, 24, 0, 28], [0, 13, 0, 17, 0, 21, 23, 0, 0, 29], [0, 14, 0, 0, 0, 22, 24, 0, 0, 30], [0, 15, 0, 0, 0, 0, 0, 0, 0, 31], [14, 16, 0, 20, 22, 0, 0, 0, 0, 32]]>
module BitSerialMatrixMultiplyState_WIDTH_10_HEIGHT_15_MATRIX___0_2_0_0_0_10_0_0_0_18___0_3_0_0_0_0_0_0_0_19___2_4_0_0_10_0_14_0_0_20___0_5_7_9_0_0_15_0_0_21___0_6_0_0_0_0_0_0_0_22___0_7_0_0_0_15_0_0_0_23___6_8_0_12_14_16_0_0_0_24___0_9_0_0_0_0_0_21_0_25___0_10_12_0_0_0_0_22_0_26___0_11_0_0_0_0_0_23_0_27___10_12_14_0_18_0_0_24_0_28___0_13_0_17_0_21_23_0_0_29___0_14_0_0_0_22_24_0_0_30___0_15_0_0_0_0_0_0_0_31___14_16_0_20_22_0_0_0_0_32___(
	input clk,
	input wire  start,
	input wire  feed,
	input wire [9:0] vector_bits,
	output /*state*/ logic [14:0][31:0] result_vector
);

/*latency*/ logic  _feed_N2; always_ff @(posedge clk) begin _feed_N2 <= feed; end
/*latency*/ logic  _feed_N1; always_ff @(posedge clk) begin _feed_N1 <= _feed_N2; end
/*latency*/ logic  _feed_D0; always_ff @(posedge clk) begin _feed_D0 <= _feed_N1; end
wire [31:0] _2 = result_vector[0];
wire [31:0] _4 = _2 * 2;
/*mux_wire*/ logic [9:0] row_bits;
wire [31:0] row_row_total;
/*latency*/ logic [31:0] _row_row_total_D0; always_ff @(posedge clk) begin _row_row_total_D0 <= row_row_total; end
wire [31:0] _5 = _4 + _row_row_total_D0;
wire [31:0] _10 = result_vector[1];
wire [31:0] _12 = _10 * 2;
/*mux_wire*/ logic [9:0] row_2_bits;
wire [31:0] row_2_row_total;
/*latency*/ logic [31:0] _row_2_row_total_N1; always_ff @(posedge clk) begin _row_2_row_total_N1 <= row_2_row_total; end
/*latency*/ logic [31:0] _row_2_row_total_D0; always_ff @(posedge clk) begin _row_2_row_total_D0 <= _row_2_row_total_N1; end
wire [31:0] _13 = _12 + _row_2_row_total_D0;
wire [31:0] _18 = result_vector[2];
wire [31:0] _20 = _18 * 2;
/*mux_wire*/ logic [9:0] row_3_bits;
wire [31:0] row_3_row_total;
wire [31:0] _21 = _20 + row_3_row_total;
wire [31:0] _26 = result_vector[3];
wire [31:0] _28 = _26 * 2;
/*mux_wire*/ logic [9:0] row_4_bits;
wire [31:0] row_4_row_total;
wire [31:0] _29 = _28 + row_4_row_total;
wire [31:0] _34 = result_vector[4];
wire [31:0] _36 = _34 * 2;
/*mux_wire*/ logic [9:0] row_5_bits;
wire [31:0] row_5_row_total;
/*latency*/ logic [31:0] _row_5_row_total_N1; always_ff @(posedge clk) begin _row_5_row_total_N1 <= row_5_row_total; end
/*latency*/ logic [31:0] _row_5_row_total_D0; always_ff @(posedge clk) begin _row_5_row_total_D0 <= _row_5_row_total_N1; end
wire [31:0] _37 = _36 + _row_5_row_total_D0;
wire [31:0] _42 = result_vector[5];
wire [31:0] _44 = _42 * 2;
/*mux_wire*/ logic [9:0] row_6_bits;
wire [31:0] row_6_row_total;
/*latency*/ logic [31:0] _row_6_row_total_D0; always_ff @(posedge clk) begin _row_6_row_total_D0 <= row_6_row_total; end
wire [31:0] _45 = _44 + _row_6_row_total_D0;
wire [31:0] _50 = result_vector[6];
wire [31:0] _52 = _50 * 2;
/*mux_wire*/ logic [9:0] row_7_bits;
wire [31:0] row_7_row_total;
wire [31:0] _53 = _52 + row_7_row_total;
wire [31:0] _58 = result_vector[7];
wire [31:0] _60 = _58 * 2;
/*mux_wire*/ logic [9:0] row_8_bits;
wire [31:0] row_8_row_total;
/*latency*/ logic [31:0] _row_8_row_total_D0; always_ff @(posedge clk) begin _row_8_row_total_D0 <= row_8_row_total; end
wire [31:0] _61 = _60 + _row_8_row_total_D0;
wire [31:0] _66 = result_vector[8];
wire [31:0] _68 = _66 * 2;
/*mux_wire*/ logic [9:0] row_9_bits;
wire [31:0] row_9_row_total;
/*latency*/ logic [31:0] _row_9_row_total_D0; always_ff @(posedge clk) begin _row_9_row_total_D0 <= row_9_row_total; end
wire [31:0] _69 = _68 + _row_9_row_total_D0;
wire [31:0] _74 = result_vector[9];
wire [31:0] _76 = _74 * 2;
/*mux_wire*/ logic [9:0] row_10_bits;
wire [31:0] row_10_row_total;
/*latency*/ logic [31:0] _row_10_row_total_D0; always_ff @(posedge clk) begin _row_10_row_total_D0 <= row_10_row_total; end
wire [31:0] _77 = _76 + _row_10_row_total_D0;
wire [31:0] _82 = result_vector[10];
wire [31:0] _84 = _82 * 2;
/*mux_wire*/ logic [9:0] row_11_bits;
wire [31:0] row_11_row_total;
wire [31:0] _85 = _84 + row_11_row_total;
wire [31:0] _90 = result_vector[11];
wire [31:0] _92 = _90 * 2;
/*mux_wire*/ logic [9:0] row_12_bits;
wire [31:0] row_12_row_total;
wire [31:0] _93 = _92 + row_12_row_total;
wire [31:0] _98 = result_vector[12];
wire [31:0] _100 = _98 * 2;
/*mux_wire*/ logic [9:0] row_13_bits;
wire [31:0] row_13_row_total;
/*latency*/ logic [31:0] _row_13_row_total_D0; always_ff @(posedge clk) begin _row_13_row_total_D0 <= row_13_row_total; end
wire [31:0] _101 = _100 + _row_13_row_total_D0;
wire [31:0] _106 = result_vector[13];
wire [31:0] _108 = _106 * 2;
/*mux_wire*/ logic [9:0] row_14_bits;
wire [31:0] row_14_row_total;
/*latency*/ logic [31:0] _row_14_row_total_N1; always_ff @(posedge clk) begin _row_14_row_total_N1 <= row_14_row_total; end
/*latency*/ logic [31:0] _row_14_row_total_D0; always_ff @(posedge clk) begin _row_14_row_total_D0 <= _row_14_row_total_N1; end
wire [31:0] _109 = _108 + _row_14_row_total_D0;
wire [31:0] _114 = result_vector[14];
wire [31:0] _116 = _114 * 2;
/*mux_wire*/ logic [9:0] row_15_bits;
wire [31:0] row_15_row_total;
wire [31:0] _117 = _116 + row_15_row_total;
BitSerialRow_SIZE_10_WEIGHTS__0_2_0_0_0_10_0_0_0_18__ row(
	.clk(clk),
	.bits(row_bits),
	.row_total(row_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_3_0_0_0_0_0_0_0_19__ row_2(
	.clk(clk),
	.bits(row_2_bits),
	.row_total(row_2_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__2_4_0_0_10_0_14_0_0_20__ row_3(
	.clk(clk),
	.bits(row_3_bits),
	.row_total(row_3_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_5_7_9_0_0_15_0_0_21__ row_4(
	.clk(clk),
	.bits(row_4_bits),
	.row_total(row_4_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_6_0_0_0_0_0_0_0_22__ row_5(
	.clk(clk),
	.bits(row_5_bits),
	.row_total(row_5_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_7_0_0_0_15_0_0_0_23__ row_6(
	.clk(clk),
	.bits(row_6_bits),
	.row_total(row_6_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__6_8_0_12_14_16_0_0_0_24__ row_7(
	.clk(clk),
	.bits(row_7_bits),
	.row_total(row_7_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_9_0_0_0_0_0_21_0_25__ row_8(
	.clk(clk),
	.bits(row_8_bits),
	.row_total(row_8_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_10_12_0_0_0_0_22_0_26__ row_9(
	.clk(clk),
	.bits(row_9_bits),
	.row_total(row_9_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_11_0_0_0_0_0_23_0_27__ row_10(
	.clk(clk),
	.bits(row_10_bits),
	.row_total(row_10_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__10_12_14_0_18_0_0_24_0_28__ row_11(
	.clk(clk),
	.bits(row_11_bits),
	.row_total(row_11_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_13_0_17_0_21_23_0_0_29__ row_12(
	.clk(clk),
	.bits(row_12_bits),
	.row_total(row_12_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_14_0_0_0_22_24_0_0_30__ row_13(
	.clk(clk),
	.bits(row_13_bits),
	.row_total(row_13_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__0_15_0_0_0_0_0_0_0_31__ row_14(
	.clk(clk),
	.bits(row_14_bits),
	.row_total(row_14_row_total)
);
BitSerialRow_SIZE_10_WEIGHTS__14_16_0_20_22_0_0_0_0_32__ row_15(
	.clk(clk),
	.bits(row_15_bits),
	.row_total(row_15_row_total)
);
always_ff @(posedge clk) begin
	if(_feed_D0) result_vector[0] <= _5;
	if(start) result_vector[0] <= 0;
	if(_feed_D0) result_vector[1] <= _13;
	if(start) result_vector[1] <= 0;
	if(_feed_D0) result_vector[2] <= _21;
	if(start) result_vector[2] <= 0;
	if(_feed_D0) result_vector[3] <= _29;
	if(start) result_vector[3] <= 0;
	if(_feed_D0) result_vector[4] <= _37;
	if(start) result_vector[4] <= 0;
	if(_feed_D0) result_vector[5] <= _45;
	if(start) result_vector[5] <= 0;
	if(_feed_D0) result_vector[6] <= _53;
	if(start) result_vector[6] <= 0;
	if(_feed_D0) result_vector[7] <= _61;
	if(start) result_vector[7] <= 0;
	if(_feed_D0) result_vector[8] <= _69;
	if(start) result_vector[8] <= 0;
	if(_feed_D0) result_vector[9] <= _77;
	if(start) result_vector[9] <= 0;
	if(_feed_D0) result_vector[10] <= _85;
	if(start) result_vector[10] <= 0;
	if(_feed_D0) result_vector[11] <= _93;
	if(start) result_vector[11] <= 0;
	if(_feed_D0) result_vector[12] <= _101;
	if(start) result_vector[12] <= 0;
	if(_feed_D0) result_vector[13] <= _109;
	if(start) result_vector[13] <= 0;
	if(_feed_D0) result_vector[14] <= _117;
	if(start) result_vector[14] <= 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_bits[0] = 'x;
	row_bits[1] = 'x;
	row_bits[2] = 'x;
	row_bits[3] = 'x;
	row_bits[4] = 'x;
	row_bits[5] = 'x;
	row_bits[6] = 'x;
	row_bits[7] = 'x;
	row_bits[8] = 'x;
	row_bits[9] = 'x;
	if(feed) row_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_2_bits[0] = 'x;
	row_2_bits[1] = 'x;
	row_2_bits[2] = 'x;
	row_2_bits[3] = 'x;
	row_2_bits[4] = 'x;
	row_2_bits[5] = 'x;
	row_2_bits[6] = 'x;
	row_2_bits[7] = 'x;
	row_2_bits[8] = 'x;
	row_2_bits[9] = 'x;
	if(feed) row_2_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_3_bits[0] = 'x;
	row_3_bits[1] = 'x;
	row_3_bits[2] = 'x;
	row_3_bits[3] = 'x;
	row_3_bits[4] = 'x;
	row_3_bits[5] = 'x;
	row_3_bits[6] = 'x;
	row_3_bits[7] = 'x;
	row_3_bits[8] = 'x;
	row_3_bits[9] = 'x;
	if(feed) row_3_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_4_bits[0] = 'x;
	row_4_bits[1] = 'x;
	row_4_bits[2] = 'x;
	row_4_bits[3] = 'x;
	row_4_bits[4] = 'x;
	row_4_bits[5] = 'x;
	row_4_bits[6] = 'x;
	row_4_bits[7] = 'x;
	row_4_bits[8] = 'x;
	row_4_bits[9] = 'x;
	if(feed) row_4_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_5_bits[0] = 'x;
	row_5_bits[1] = 'x;
	row_5_bits[2] = 'x;
	row_5_bits[3] = 'x;
	row_5_bits[4] = 'x;
	row_5_bits[5] = 'x;
	row_5_bits[6] = 'x;
	row_5_bits[7] = 'x;
	row_5_bits[8] = 'x;
	row_5_bits[9] = 'x;
	if(feed) row_5_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_6_bits[0] = 'x;
	row_6_bits[1] = 'x;
	row_6_bits[2] = 'x;
	row_6_bits[3] = 'x;
	row_6_bits[4] = 'x;
	row_6_bits[5] = 'x;
	row_6_bits[6] = 'x;
	row_6_bits[7] = 'x;
	row_6_bits[8] = 'x;
	row_6_bits[9] = 'x;
	if(feed) row_6_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_7_bits[0] = 'x;
	row_7_bits[1] = 'x;
	row_7_bits[2] = 'x;
	row_7_bits[3] = 'x;
	row_7_bits[4] = 'x;
	row_7_bits[5] = 'x;
	row_7_bits[6] = 'x;
	row_7_bits[7] = 'x;
	row_7_bits[8] = 'x;
	row_7_bits[9] = 'x;
	if(feed) row_7_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_8_bits[0] = 'x;
	row_8_bits[1] = 'x;
	row_8_bits[2] = 'x;
	row_8_bits[3] = 'x;
	row_8_bits[4] = 'x;
	row_8_bits[5] = 'x;
	row_8_bits[6] = 'x;
	row_8_bits[7] = 'x;
	row_8_bits[8] = 'x;
	row_8_bits[9] = 'x;
	if(feed) row_8_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_9_bits[0] = 'x;
	row_9_bits[1] = 'x;
	row_9_bits[2] = 'x;
	row_9_bits[3] = 'x;
	row_9_bits[4] = 'x;
	row_9_bits[5] = 'x;
	row_9_bits[6] = 'x;
	row_9_bits[7] = 'x;
	row_9_bits[8] = 'x;
	row_9_bits[9] = 'x;
	if(feed) row_9_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_10_bits[0] = 'x;
	row_10_bits[1] = 'x;
	row_10_bits[2] = 'x;
	row_10_bits[3] = 'x;
	row_10_bits[4] = 'x;
	row_10_bits[5] = 'x;
	row_10_bits[6] = 'x;
	row_10_bits[7] = 'x;
	row_10_bits[8] = 'x;
	row_10_bits[9] = 'x;
	if(feed) row_10_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_11_bits[0] = 'x;
	row_11_bits[1] = 'x;
	row_11_bits[2] = 'x;
	row_11_bits[3] = 'x;
	row_11_bits[4] = 'x;
	row_11_bits[5] = 'x;
	row_11_bits[6] = 'x;
	row_11_bits[7] = 'x;
	row_11_bits[8] = 'x;
	row_11_bits[9] = 'x;
	if(feed) row_11_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_12_bits[0] = 'x;
	row_12_bits[1] = 'x;
	row_12_bits[2] = 'x;
	row_12_bits[3] = 'x;
	row_12_bits[4] = 'x;
	row_12_bits[5] = 'x;
	row_12_bits[6] = 'x;
	row_12_bits[7] = 'x;
	row_12_bits[8] = 'x;
	row_12_bits[9] = 'x;
	if(feed) row_12_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_13_bits[0] = 'x;
	row_13_bits[1] = 'x;
	row_13_bits[2] = 'x;
	row_13_bits[3] = 'x;
	row_13_bits[4] = 'x;
	row_13_bits[5] = 'x;
	row_13_bits[6] = 'x;
	row_13_bits[7] = 'x;
	row_13_bits[8] = 'x;
	row_13_bits[9] = 'x;
	if(feed) row_13_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_14_bits[0] = 'x;
	row_14_bits[1] = 'x;
	row_14_bits[2] = 'x;
	row_14_bits[3] = 'x;
	row_14_bits[4] = 'x;
	row_14_bits[5] = 'x;
	row_14_bits[6] = 'x;
	row_14_bits[7] = 'x;
	row_14_bits[8] = 'x;
	row_14_bits[9] = 'x;
	if(feed) row_14_bits = vector_bits;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_15_bits[0] = 'x;
	row_15_bits[1] = 'x;
	row_15_bits[2] = 'x;
	row_15_bits[3] = 'x;
	row_15_bits[4] = 'x;
	row_15_bits[5] = 'x;
	row_15_bits[6] = 'x;
	row_15_bits[7] = 'x;
	row_15_bits[8] = 'x;
	row_15_bits[9] = 'x;
	if(feed) row_15_bits = vector_bits;
end
endmodule

// ::FixedSizeIterator::<UP_TO = 32>
module FixedSizeIterator_UP_TO_32_(
	input clk,
	output /*mux_wire*/ logic  valid,
	output /*state*/ logic [31:0] value,
	output /*mux_wire*/ logic  last,
	input wire  start
);

wire  _2 = value == 31;
wire  _4 = value != 32;
wire [31:0] _7 = value + 1;
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	valid = 'x;
	valid = _4;
end
always_ff @(posedge clk) begin
	if(start) value <= 0;
	if(!start) if(valid) value <= _7;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	last = 'x;
	last = _2;
end
endmodule

// ::LatencyOffset::<T = ::int[15], OFFSET = 33>
module LatencyOffset_T_int_15__OFFSET_33_(
	input clk,
	input wire [14:0][31:0] in,
	output /*mux_wire*/ logic [14:0][31:0] out
);

	assign out = in;
endmodule

// ::IntToBits
module IntToBits(
	input clk,
	input wire [31:0] value,
	output /*mux_wire*/ logic [31:0] bits
);

	assign bits[0] = value[0];
	assign bits[1] = value[1];
	assign bits[2] = value[2];
	assign bits[3] = value[3];
	assign bits[4] = value[4];
	assign bits[5] = value[5];
	assign bits[6] = value[6];
	assign bits[7] = value[7];
	assign bits[8] = value[8];
	assign bits[9] = value[9];
	assign bits[10] = value[10];
	assign bits[11] = value[11];
	assign bits[12] = value[12];
	assign bits[13] = value[13];
	assign bits[14] = value[14];
	assign bits[15] = value[15];
	assign bits[16] = value[16];
	assign bits[17] = value[17];
	assign bits[18] = value[18];
	assign bits[19] = value[19];
	assign bits[20] = value[20];
	assign bits[21] = value[21];
	assign bits[22] = value[22];
	assign bits[23] = value[23];
	assign bits[24] = value[24];
	assign bits[25] = value[25];
	assign bits[26] = value[26];
	assign bits[27] = value[27];
	assign bits[28] = value[28];
	assign bits[29] = value[29];
	assign bits[30] = value[30];
	assign bits[31] = value[31];
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 2, 0, 0, 0, 10, 0, 0, 0, 18]>
module BitSerialRow_SIZE_10_WEIGHTS__0_2_0_0_0_10_0_0_0_18__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [2:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[5];
wire  _14 = bits[9];
/*mux_wire*/ logic [2:0][31:0] _19_values;
wire [31:0] _19_total;
TreeAdd_WIDTH_3_ _19(
	.clk(clk),
	.values(_19_values),
	.total(_19_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _19_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	if(_2) nonzero_weights[0] = 2;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 10;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 18;
	if(!_14) nonzero_weights[2] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_19_values[0] = 'x;
	_19_values[1] = 'x;
	_19_values[2] = 'x;
	_19_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 3, 0, 0, 0, 0, 0, 0, 0, 19]>
module BitSerialRow_SIZE_10_WEIGHTS__0_3_0_0_0_0_0_0_0_19__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [1:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[9];
/*mux_wire*/ logic [1:0][31:0] _13_values;
wire [31:0] _13_total;
TreeAdd_WIDTH_2_ _13(
	.clk(clk),
	.values(_13_values),
	.total(_13_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _13_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	if(_2) nonzero_weights[0] = 3;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 19;
	if(!_8) nonzero_weights[1] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_13_values[0] = 'x;
	_13_values[1] = 'x;
	_13_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [2, 4, 0, 0, 10, 0, 14, 0, 0, 20]>
module BitSerialRow_SIZE_10_WEIGHTS__2_4_0_0_10_0_14_0_0_20__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [4:0][31:0] nonzero_weights;
wire  _2 = bits[0];
wire  _8 = bits[1];
wire  _14 = bits[4];
wire  _20 = bits[6];
wire  _26 = bits[9];
/*mux_wire*/ logic [4:0][31:0] _31_values;
wire [31:0] _31_total;
TreeAdd_WIDTH_5_ _31(
	.clk(clk),
	.values(_31_values),
	.total(_31_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _31_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	nonzero_weights[4] = 'x;
	if(_2) nonzero_weights[0] = 2;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 4;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 10;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 14;
	if(!_20) nonzero_weights[3] = 0;
	if(_26) nonzero_weights[4] = 20;
	if(!_26) nonzero_weights[4] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_31_values[0] = 'x;
	_31_values[1] = 'x;
	_31_values[2] = 'x;
	_31_values[3] = 'x;
	_31_values[4] = 'x;
	_31_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 5, 7, 9, 0, 0, 15, 0, 0, 21]>
module BitSerialRow_SIZE_10_WEIGHTS__0_5_7_9_0_0_15_0_0_21__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [4:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[2];
wire  _14 = bits[3];
wire  _20 = bits[6];
wire  _26 = bits[9];
/*mux_wire*/ logic [4:0][31:0] _31_values;
wire [31:0] _31_total;
TreeAdd_WIDTH_5_ _31(
	.clk(clk),
	.values(_31_values),
	.total(_31_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _31_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	nonzero_weights[4] = 'x;
	if(_2) nonzero_weights[0] = 5;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 7;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 9;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 15;
	if(!_20) nonzero_weights[3] = 0;
	if(_26) nonzero_weights[4] = 21;
	if(!_26) nonzero_weights[4] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_31_values[0] = 'x;
	_31_values[1] = 'x;
	_31_values[2] = 'x;
	_31_values[3] = 'x;
	_31_values[4] = 'x;
	_31_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 6, 0, 0, 0, 0, 0, 0, 0, 22]>
module BitSerialRow_SIZE_10_WEIGHTS__0_6_0_0_0_0_0_0_0_22__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [1:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[9];
/*mux_wire*/ logic [1:0][31:0] _13_values;
wire [31:0] _13_total;
TreeAdd_WIDTH_2_ _13(
	.clk(clk),
	.values(_13_values),
	.total(_13_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _13_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	if(_2) nonzero_weights[0] = 6;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 22;
	if(!_8) nonzero_weights[1] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_13_values[0] = 'x;
	_13_values[1] = 'x;
	_13_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 7, 0, 0, 0, 15, 0, 0, 0, 23]>
module BitSerialRow_SIZE_10_WEIGHTS__0_7_0_0_0_15_0_0_0_23__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [2:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[5];
wire  _14 = bits[9];
/*mux_wire*/ logic [2:0][31:0] _19_values;
wire [31:0] _19_total;
TreeAdd_WIDTH_3_ _19(
	.clk(clk),
	.values(_19_values),
	.total(_19_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _19_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	if(_2) nonzero_weights[0] = 7;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 15;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 23;
	if(!_14) nonzero_weights[2] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_19_values[0] = 'x;
	_19_values[1] = 'x;
	_19_values[2] = 'x;
	_19_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [6, 8, 0, 12, 14, 16, 0, 0, 0, 24]>
module BitSerialRow_SIZE_10_WEIGHTS__6_8_0_12_14_16_0_0_0_24__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [5:0][31:0] nonzero_weights;
wire  _2 = bits[0];
wire  _8 = bits[1];
wire  _14 = bits[3];
wire  _20 = bits[4];
wire  _26 = bits[5];
wire  _32 = bits[9];
/*mux_wire*/ logic [5:0][31:0] _37_values;
wire [31:0] _37_total;
TreeAdd_WIDTH_6_ _37(
	.clk(clk),
	.values(_37_values),
	.total(_37_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _37_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	nonzero_weights[4] = 'x;
	nonzero_weights[5] = 'x;
	if(_2) nonzero_weights[0] = 6;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 8;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 12;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 14;
	if(!_20) nonzero_weights[3] = 0;
	if(_26) nonzero_weights[4] = 16;
	if(!_26) nonzero_weights[4] = 0;
	if(_32) nonzero_weights[5] = 24;
	if(!_32) nonzero_weights[5] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_37_values[0] = 'x;
	_37_values[1] = 'x;
	_37_values[2] = 'x;
	_37_values[3] = 'x;
	_37_values[4] = 'x;
	_37_values[5] = 'x;
	_37_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 9, 0, 0, 0, 0, 0, 21, 0, 25]>
module BitSerialRow_SIZE_10_WEIGHTS__0_9_0_0_0_0_0_21_0_25__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [2:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[7];
wire  _14 = bits[9];
/*mux_wire*/ logic [2:0][31:0] _19_values;
wire [31:0] _19_total;
TreeAdd_WIDTH_3_ _19(
	.clk(clk),
	.values(_19_values),
	.total(_19_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _19_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	if(_2) nonzero_weights[0] = 9;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 21;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 25;
	if(!_14) nonzero_weights[2] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_19_values[0] = 'x;
	_19_values[1] = 'x;
	_19_values[2] = 'x;
	_19_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 10, 12, 0, 0, 0, 0, 22, 0, 26]>
module BitSerialRow_SIZE_10_WEIGHTS__0_10_12_0_0_0_0_22_0_26__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [3:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[2];
wire  _14 = bits[7];
wire  _20 = bits[9];
/*mux_wire*/ logic [3:0][31:0] _25_values;
wire [31:0] _25_total;
TreeAdd_WIDTH_4_ _25(
	.clk(clk),
	.values(_25_values),
	.total(_25_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _25_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	if(_2) nonzero_weights[0] = 10;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 12;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 22;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 26;
	if(!_20) nonzero_weights[3] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_25_values[0] = 'x;
	_25_values[1] = 'x;
	_25_values[2] = 'x;
	_25_values[3] = 'x;
	_25_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 11, 0, 0, 0, 0, 0, 23, 0, 27]>
module BitSerialRow_SIZE_10_WEIGHTS__0_11_0_0_0_0_0_23_0_27__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [2:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[7];
wire  _14 = bits[9];
/*mux_wire*/ logic [2:0][31:0] _19_values;
wire [31:0] _19_total;
TreeAdd_WIDTH_3_ _19(
	.clk(clk),
	.values(_19_values),
	.total(_19_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _19_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	if(_2) nonzero_weights[0] = 11;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 23;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 27;
	if(!_14) nonzero_weights[2] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_19_values[0] = 'x;
	_19_values[1] = 'x;
	_19_values[2] = 'x;
	_19_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [10, 12, 14, 0, 18, 0, 0, 24, 0, 28]>
module BitSerialRow_SIZE_10_WEIGHTS__10_12_14_0_18_0_0_24_0_28__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [5:0][31:0] nonzero_weights;
wire  _2 = bits[0];
wire  _8 = bits[1];
wire  _14 = bits[2];
wire  _20 = bits[4];
wire  _26 = bits[7];
wire  _32 = bits[9];
/*mux_wire*/ logic [5:0][31:0] _37_values;
wire [31:0] _37_total;
TreeAdd_WIDTH_6_ _37(
	.clk(clk),
	.values(_37_values),
	.total(_37_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _37_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	nonzero_weights[4] = 'x;
	nonzero_weights[5] = 'x;
	if(_2) nonzero_weights[0] = 10;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 12;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 14;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 18;
	if(!_20) nonzero_weights[3] = 0;
	if(_26) nonzero_weights[4] = 24;
	if(!_26) nonzero_weights[4] = 0;
	if(_32) nonzero_weights[5] = 28;
	if(!_32) nonzero_weights[5] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_37_values[0] = 'x;
	_37_values[1] = 'x;
	_37_values[2] = 'x;
	_37_values[3] = 'x;
	_37_values[4] = 'x;
	_37_values[5] = 'x;
	_37_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 13, 0, 17, 0, 21, 23, 0, 0, 29]>
module BitSerialRow_SIZE_10_WEIGHTS__0_13_0_17_0_21_23_0_0_29__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [4:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[3];
wire  _14 = bits[5];
wire  _20 = bits[6];
wire  _26 = bits[9];
/*mux_wire*/ logic [4:0][31:0] _31_values;
wire [31:0] _31_total;
TreeAdd_WIDTH_5_ _31(
	.clk(clk),
	.values(_31_values),
	.total(_31_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _31_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	nonzero_weights[4] = 'x;
	if(_2) nonzero_weights[0] = 13;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 17;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 21;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 23;
	if(!_20) nonzero_weights[3] = 0;
	if(_26) nonzero_weights[4] = 29;
	if(!_26) nonzero_weights[4] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_31_values[0] = 'x;
	_31_values[1] = 'x;
	_31_values[2] = 'x;
	_31_values[3] = 'x;
	_31_values[4] = 'x;
	_31_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 14, 0, 0, 0, 22, 24, 0, 0, 30]>
module BitSerialRow_SIZE_10_WEIGHTS__0_14_0_0_0_22_24_0_0_30__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [3:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[5];
wire  _14 = bits[6];
wire  _20 = bits[9];
/*mux_wire*/ logic [3:0][31:0] _25_values;
wire [31:0] _25_total;
TreeAdd_WIDTH_4_ _25(
	.clk(clk),
	.values(_25_values),
	.total(_25_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _25_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	if(_2) nonzero_weights[0] = 14;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 22;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 24;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 30;
	if(!_20) nonzero_weights[3] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_25_values[0] = 'x;
	_25_values[1] = 'x;
	_25_values[2] = 'x;
	_25_values[3] = 'x;
	_25_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [0, 15, 0, 0, 0, 0, 0, 0, 0, 31]>
module BitSerialRow_SIZE_10_WEIGHTS__0_15_0_0_0_0_0_0_0_31__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [1:0][31:0] nonzero_weights;
wire  _2 = bits[1];
wire  _8 = bits[9];
/*mux_wire*/ logic [1:0][31:0] _13_values;
wire [31:0] _13_total;
TreeAdd_WIDTH_2_ _13(
	.clk(clk),
	.values(_13_values),
	.total(_13_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _13_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	if(_2) nonzero_weights[0] = 15;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 31;
	if(!_8) nonzero_weights[1] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_13_values[0] = 'x;
	_13_values[1] = 'x;
	_13_values = nonzero_weights;
end
endmodule

// ::BitSerialRow::<SIZE = 10, WEIGHTS = [14, 16, 0, 20, 22, 0, 0, 0, 0, 32]>
module BitSerialRow_SIZE_10_WEIGHTS__14_16_0_20_22_0_0_0_0_32__(
	input clk,
	input wire [9:0] bits,
	output /*mux_wire*/ logic [31:0] row_total
);

/*mux_wire*/ logic [4:0][31:0] nonzero_weights;
wire  _2 = bits[0];
wire  _8 = bits[1];
wire  _14 = bits[3];
wire  _20 = bits[4];
wire  _26 = bits[9];
/*mux_wire*/ logic [4:0][31:0] _31_values;
wire [31:0] _31_total;
TreeAdd_WIDTH_5_ _31(
	.clk(clk),
	.values(_31_values),
	.total(_31_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	row_total = 'x;
	row_total = _31_total;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	nonzero_weights[0] = 'x;
	nonzero_weights[1] = 'x;
	nonzero_weights[2] = 'x;
	nonzero_weights[3] = 'x;
	nonzero_weights[4] = 'x;
	if(_2) nonzero_weights[0] = 14;
	if(!_2) nonzero_weights[0] = 0;
	if(_8) nonzero_weights[1] = 16;
	if(!_8) nonzero_weights[1] = 0;
	if(_14) nonzero_weights[2] = 20;
	if(!_14) nonzero_weights[2] = 0;
	if(_20) nonzero_weights[3] = 22;
	if(!_20) nonzero_weights[3] = 0;
	if(_26) nonzero_weights[4] = 32;
	if(!_26) nonzero_weights[4] = 0;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_31_values[0] = 'x;
	_31_values[1] = 'x;
	_31_values[2] = 'x;
	_31_values[3] = 'x;
	_31_values[4] = 'x;
	_31_values = nonzero_weights;
end
endmodule

// ::TreeAdd::<WIDTH = 3>
module TreeAdd_WIDTH_3_(
	input clk,
	input wire [2:0][31:0] values,
	output /*mux_wire*/ logic [31:0] total
);

/*mux_wire*/ logic [0:0][31:0] left_part;
/*mux_wire*/ logic [1:0][31:0] right_part;
/*mux_wire*/ logic [2:0][31:0] _1_i;
wire [0:0][31:0] _1_left;
wire [1:0][31:0] _1_right;
/*mux_wire*/ logic [0:0][31:0] _2_values;
wire [31:0] _2_total;
/*latency*/ logic [31:0] __2_total_D1; always_ff @(posedge clk) begin __2_total_D1 <= _2_total; end
/*mux_wire*/ logic [1:0][31:0] _3_values;
wire [31:0] _3_total;
wire [31:0] _4 = __2_total_D1 + _3_total;
/*latency*/ logic [31:0] __4_D2; always_ff @(posedge clk) begin __4_D2 <= _4; end
SplitAt_T_int_SIZE_3_SPLIT_POINT_1_ _1(
	.clk(clk),
	.i(_1_i),
	.left(_1_left),
	.right(_1_right)
);
TreeAdd_WIDTH_1_ _2(
	.clk(clk),
	.values(_2_values),
	.total(_2_total)
);
TreeAdd_WIDTH_2_ _3(
	.clk(clk),
	.values(_3_values),
	.total(_3_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	total = 'x;
	total = __4_D2;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left_part[0] = 'x;
	left_part = _1_left;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right_part[0] = 'x;
	right_part[1] = 'x;
	right_part = _1_right;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1_i[0] = 'x;
	_1_i[1] = 'x;
	_1_i[2] = 'x;
	_1_i = values;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_2_values[0] = 'x;
	_2_values = left_part;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_3_values[0] = 'x;
	_3_values[1] = 'x;
	_3_values = right_part;
end
endmodule

// ::TreeAdd::<WIDTH = 2>
module TreeAdd_WIDTH_2_(
	input clk,
	input wire [1:0][31:0] values,
	output /*mux_wire*/ logic [31:0] total
);

/*mux_wire*/ logic [0:0][31:0] left_part;
/*mux_wire*/ logic [0:0][31:0] right_part;
/*mux_wire*/ logic [1:0][31:0] _1_i;
wire [0:0][31:0] _1_left;
wire [0:0][31:0] _1_right;
/*mux_wire*/ logic [0:0][31:0] _2_values;
wire [31:0] _2_total;
/*mux_wire*/ logic [0:0][31:0] _3_values;
wire [31:0] _3_total;
wire [31:0] _4 = _2_total + _3_total;
/*latency*/ logic [31:0] __4_D1; always_ff @(posedge clk) begin __4_D1 <= _4; end
SplitAt_T_int_SIZE_2_SPLIT_POINT_1_ _1(
	.clk(clk),
	.i(_1_i),
	.left(_1_left),
	.right(_1_right)
);
TreeAdd_WIDTH_1_ _2(
	.clk(clk),
	.values(_2_values),
	.total(_2_total)
);
TreeAdd_WIDTH_1_ _3(
	.clk(clk),
	.values(_3_values),
	.total(_3_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	total = 'x;
	total = __4_D1;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left_part[0] = 'x;
	left_part = _1_left;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right_part[0] = 'x;
	right_part = _1_right;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1_i[0] = 'x;
	_1_i[1] = 'x;
	_1_i = values;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_2_values[0] = 'x;
	_2_values = left_part;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_3_values[0] = 'x;
	_3_values = right_part;
end
endmodule

// ::TreeAdd::<WIDTH = 5>
module TreeAdd_WIDTH_5_(
	input clk,
	input wire [4:0][31:0] values,
	output /*mux_wire*/ logic [31:0] total
);

/*mux_wire*/ logic [1:0][31:0] left_part;
/*mux_wire*/ logic [2:0][31:0] right_part;
/*mux_wire*/ logic [4:0][31:0] _1_i;
wire [1:0][31:0] _1_left;
wire [2:0][31:0] _1_right;
/*mux_wire*/ logic [1:0][31:0] _2_values;
wire [31:0] _2_total;
/*latency*/ logic [31:0] __2_total_D2; always_ff @(posedge clk) begin __2_total_D2 <= _2_total; end
/*mux_wire*/ logic [2:0][31:0] _3_values;
wire [31:0] _3_total;
wire [31:0] _4 = __2_total_D2 + _3_total;
/*latency*/ logic [31:0] __4_D3; always_ff @(posedge clk) begin __4_D3 <= _4; end
SplitAt_T_int_SIZE_5_SPLIT_POINT_2_ _1(
	.clk(clk),
	.i(_1_i),
	.left(_1_left),
	.right(_1_right)
);
TreeAdd_WIDTH_2_ _2(
	.clk(clk),
	.values(_2_values),
	.total(_2_total)
);
TreeAdd_WIDTH_3_ _3(
	.clk(clk),
	.values(_3_values),
	.total(_3_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	total = 'x;
	total = __4_D3;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left_part[0] = 'x;
	left_part[1] = 'x;
	left_part = _1_left;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right_part[0] = 'x;
	right_part[1] = 'x;
	right_part[2] = 'x;
	right_part = _1_right;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1_i[0] = 'x;
	_1_i[1] = 'x;
	_1_i[2] = 'x;
	_1_i[3] = 'x;
	_1_i[4] = 'x;
	_1_i = values;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_2_values[0] = 'x;
	_2_values[1] = 'x;
	_2_values = left_part;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_3_values[0] = 'x;
	_3_values[1] = 'x;
	_3_values[2] = 'x;
	_3_values = right_part;
end
endmodule

// ::TreeAdd::<WIDTH = 6>
module TreeAdd_WIDTH_6_(
	input clk,
	input wire [5:0][31:0] values,
	output /*mux_wire*/ logic [31:0] total
);

/*mux_wire*/ logic [2:0][31:0] left_part;
/*mux_wire*/ logic [2:0][31:0] right_part;
/*mux_wire*/ logic [5:0][31:0] _1_i;
wire [2:0][31:0] _1_left;
wire [2:0][31:0] _1_right;
/*mux_wire*/ logic [2:0][31:0] _2_values;
wire [31:0] _2_total;
/*mux_wire*/ logic [2:0][31:0] _3_values;
wire [31:0] _3_total;
wire [31:0] _4 = _2_total + _3_total;
/*latency*/ logic [31:0] __4_D3; always_ff @(posedge clk) begin __4_D3 <= _4; end
SplitAt_T_int_SIZE_6_SPLIT_POINT_3_ _1(
	.clk(clk),
	.i(_1_i),
	.left(_1_left),
	.right(_1_right)
);
TreeAdd_WIDTH_3_ _2(
	.clk(clk),
	.values(_2_values),
	.total(_2_total)
);
TreeAdd_WIDTH_3_ _3(
	.clk(clk),
	.values(_3_values),
	.total(_3_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	total = 'x;
	total = __4_D3;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left_part[0] = 'x;
	left_part[1] = 'x;
	left_part[2] = 'x;
	left_part = _1_left;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right_part[0] = 'x;
	right_part[1] = 'x;
	right_part[2] = 'x;
	right_part = _1_right;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1_i[0] = 'x;
	_1_i[1] = 'x;
	_1_i[2] = 'x;
	_1_i[3] = 'x;
	_1_i[4] = 'x;
	_1_i[5] = 'x;
	_1_i = values;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_2_values[0] = 'x;
	_2_values[1] = 'x;
	_2_values[2] = 'x;
	_2_values = left_part;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_3_values[0] = 'x;
	_3_values[1] = 'x;
	_3_values[2] = 'x;
	_3_values = right_part;
end
endmodule

// ::TreeAdd::<WIDTH = 4>
module TreeAdd_WIDTH_4_(
	input clk,
	input wire [3:0][31:0] values,
	output /*mux_wire*/ logic [31:0] total
);

/*mux_wire*/ logic [1:0][31:0] left_part;
/*mux_wire*/ logic [1:0][31:0] right_part;
/*mux_wire*/ logic [3:0][31:0] _1_i;
wire [1:0][31:0] _1_left;
wire [1:0][31:0] _1_right;
/*mux_wire*/ logic [1:0][31:0] _2_values;
wire [31:0] _2_total;
/*mux_wire*/ logic [1:0][31:0] _3_values;
wire [31:0] _3_total;
wire [31:0] _4 = _2_total + _3_total;
/*latency*/ logic [31:0] __4_D2; always_ff @(posedge clk) begin __4_D2 <= _4; end
SplitAt_T_int_SIZE_4_SPLIT_POINT_2_ _1(
	.clk(clk),
	.i(_1_i),
	.left(_1_left),
	.right(_1_right)
);
TreeAdd_WIDTH_2_ _2(
	.clk(clk),
	.values(_2_values),
	.total(_2_total)
);
TreeAdd_WIDTH_2_ _3(
	.clk(clk),
	.values(_3_values),
	.total(_3_total)
);
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	total = 'x;
	total = __4_D2;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left_part[0] = 'x;
	left_part[1] = 'x;
	left_part = _1_left;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right_part[0] = 'x;
	right_part[1] = 'x;
	right_part = _1_right;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_1_i[0] = 'x;
	_1_i[1] = 'x;
	_1_i[2] = 'x;
	_1_i[3] = 'x;
	_1_i = values;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_2_values[0] = 'x;
	_2_values[1] = 'x;
	_2_values = left_part;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	_3_values[0] = 'x;
	_3_values[1] = 'x;
	_3_values = right_part;
end
endmodule

// ::SplitAt::<T = ::int, SIZE = 3, SPLIT_POINT = 1>
module SplitAt_T_int_SIZE_3_SPLIT_POINT_1_(
	input clk,
	input wire [2:0][31:0] i,
	output /*mux_wire*/ logic [0:0][31:0] left,
	output /*mux_wire*/ logic [1:0][31:0] right
);

wire [31:0] _2 = i[0];
wire [31:0] _5 = i[1];
wire [31:0] _8 = i[2];
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left[0] = 'x;
	left[0] = _2;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right[0] = 'x;
	right[1] = 'x;
	right[0] = _5;
	right[1] = _8;
end
endmodule

// ::TreeAdd::<WIDTH = 1>
module TreeAdd_WIDTH_1_(
	input clk,
	input wire [0:0][31:0] values,
	output /*mux_wire*/ logic [31:0] total
);

wire [31:0] _2 = values[0];
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	total = 'x;
	total = _2;
end
endmodule

// ::SplitAt::<T = ::int, SIZE = 2, SPLIT_POINT = 1>
module SplitAt_T_int_SIZE_2_SPLIT_POINT_1_(
	input clk,
	input wire [1:0][31:0] i,
	output /*mux_wire*/ logic [0:0][31:0] left,
	output /*mux_wire*/ logic [0:0][31:0] right
);

wire [31:0] _2 = i[0];
wire [31:0] _5 = i[1];
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left[0] = 'x;
	left[0] = _2;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right[0] = 'x;
	right[0] = _5;
end
endmodule

// ::SplitAt::<T = ::int, SIZE = 5, SPLIT_POINT = 2>
module SplitAt_T_int_SIZE_5_SPLIT_POINT_2_(
	input clk,
	input wire [4:0][31:0] i,
	output /*mux_wire*/ logic [1:0][31:0] left,
	output /*mux_wire*/ logic [2:0][31:0] right
);

wire [31:0] _2 = i[0];
wire [31:0] _5 = i[1];
wire [31:0] _8 = i[2];
wire [31:0] _11 = i[3];
wire [31:0] _14 = i[4];
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left[0] = 'x;
	left[1] = 'x;
	left[0] = _2;
	left[1] = _5;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right[0] = 'x;
	right[1] = 'x;
	right[2] = 'x;
	right[0] = _8;
	right[1] = _11;
	right[2] = _14;
end
endmodule

// ::SplitAt::<T = ::int, SIZE = 6, SPLIT_POINT = 3>
module SplitAt_T_int_SIZE_6_SPLIT_POINT_3_(
	input clk,
	input wire [5:0][31:0] i,
	output /*mux_wire*/ logic [2:0][31:0] left,
	output /*mux_wire*/ logic [2:0][31:0] right
);

wire [31:0] _2 = i[0];
wire [31:0] _5 = i[1];
wire [31:0] _8 = i[2];
wire [31:0] _11 = i[3];
wire [31:0] _14 = i[4];
wire [31:0] _17 = i[5];
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left[0] = 'x;
	left[1] = 'x;
	left[2] = 'x;
	left[0] = _2;
	left[1] = _5;
	left[2] = _8;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right[0] = 'x;
	right[1] = 'x;
	right[2] = 'x;
	right[0] = _11;
	right[1] = _14;
	right[2] = _17;
end
endmodule

// ::SplitAt::<T = ::int, SIZE = 4, SPLIT_POINT = 2>
module SplitAt_T_int_SIZE_4_SPLIT_POINT_2_(
	input clk,
	input wire [3:0][31:0] i,
	output /*mux_wire*/ logic [1:0][31:0] left,
	output /*mux_wire*/ logic [1:0][31:0] right
);

wire [31:0] _2 = i[0];
wire [31:0] _5 = i[1];
wire [31:0] _8 = i[2];
wire [31:0] _11 = i[3];
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	left[0] = 'x;
	left[1] = 'x;
	left[0] = _2;
	left[1] = _5;
end
always_comb begin
	// Combinatorial wires are not defined when not valid. This is just so that the synthesys tool doesn't generate latches
	right[0] = 'x;
	right[1] = 'x;
	right[0] = _8;
	right[1] = _11;
end
endmodule

